// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.0.396.4
// Netlist written on Thu Aug 13 13:06:25 2020
//
// Verilog Description of module mcm_top
//

module mcm_top (clk_in, resetn, led_sw, cs, intrpt_out, FLASH_CS, 
            MAX3421_CS, CS_READY, spi_clk, spi_mosi, spi_miso, spi_scsn, 
            UC_TXD0, UC_RXD0, pin_io, C_1, C_2, C_3, C_4, C_5, 
            C_6, C_7, C_8) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(9[8:15])
    input clk_in;   // c:/s_links/sources/mcm_top.v(16[27:33])
    input resetn;   // c:/s_links/sources/mcm_top.v(17[27:33])
    output led_sw;   // c:/s_links/sources/mcm_top.v(18[24:30])
    input [4:0]cs;   // c:/s_links/sources/mcm_top.v(19[37:39])
    output [6:0]intrpt_out;   // c:/s_links/sources/mcm_top.v(20[36:46])
    output FLASH_CS;   // c:/s_links/sources/mcm_top.v(21[24:32])
    output MAX3421_CS;   // c:/s_links/sources/mcm_top.v(22[24:34])
    input CS_READY;   // c:/s_links/sources/mcm_top.v(23[24:32])
    input spi_clk /* synthesis black_box_pad_pin=1 */ ;   // c:/s_links/sources/mcm_top.v(26[27:34])
    input spi_mosi /* synthesis black_box_pad_pin=1 */ ;   // c:/s_links/sources/mcm_top.v(27[27:35])
    output spi_miso /* synthesis black_box_pad_pin=1 */ ;   // c:/s_links/sources/mcm_top.v(28[27:35])
    input spi_scsn;   // c:/s_links/sources/mcm_top.v(29[27:35])
    input UC_TXD0;   // c:/s_links/sources/mcm_top.v(32[27:34])
    output UC_RXD0;   // c:/s_links/sources/mcm_top.v(33[27:34])
    inout [69:0]pin_io;   // c:/s_links/sources/mcm_top.v(36[51:57])
    input C_1 /* synthesis .original_dir=IN_OUT */ ;   // c:/s_links/sources/mcm_top.v(39[24:27])
    input C_2 /* synthesis .original_dir=IN_OUT */ ;   // c:/s_links/sources/mcm_top.v(40[24:27])
    input C_3 /* synthesis .original_dir=IN_OUT */ ;   // c:/s_links/sources/mcm_top.v(41[24:27])
    input C_4 /* synthesis .original_dir=IN_OUT */ ;   // c:/s_links/sources/mcm_top.v(42[24:27])
    input C_5 /* synthesis .original_dir=IN_OUT */ ;   // c:/s_links/sources/mcm_top.v(43[24:27])
    input C_6 /* synthesis .original_dir=IN_OUT */ ;   // c:/s_links/sources/mcm_top.v(44[24:27])
    output C_7 /* synthesis .original_dir=IN_OUT */ ;   // c:/s_links/sources/mcm_top.v(45[24:27])
    input C_8 /* synthesis .original_dir=IN_OUT */ ;   // c:/s_links/sources/mcm_top.v(46[24:27])
    
    wire clk_in_c /* synthesis is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(16[27:33])
    wire CS_READY_c /* synthesis is_clock=1, SET_AS_NETWORK=CS_READY_c */ ;   // c:/s_links/sources/mcm_top.v(23[24:32])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire [20:0]pin_intrpt /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[20] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    wire clk_100k /* synthesis SET_AS_NETWORK=clk_100k, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(134[6:14])
    wire clk_1MHz /* synthesis SET_AS_NETWORK=clk_1MHz, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(136[6:14])
    wire spi_clk_i /* synthesis is_clock=1 */ ;   // c:/s_links/sources/config_hex/ip/spi_slave_efb.v(34[10:19])
    
    wire GND_net, resetn_c, led_sw_c, cs_c_4, cs_c_3, cs_c_2, cs_c_1, 
        cs_c_0, intrpt_out_c_6, intrpt_out_c_5, intrpt_out_c_4, intrpt_out_c_3, 
        intrpt_out_c_2, intrpt_out_c_1, intrpt_out_c_0, FLASH_CS_c, 
        MAX3421_CS_c, spi_scsn_c, UC_TXD0_c, pin_io_c_68, pin_io_c_64, 
        pin_io_c_63, pin_io_c_62, pin_io_c_58, pin_io_c_54, pin_io_c_53, 
        pin_io_c_52, pin_io_c_48, pin_io_c_44, pin_io_c_43, pin_io_c_42, 
        pin_io_c_38, pin_io_c_34, pin_io_c_33, pin_io_c_32, pin_io_c_28, 
        pin_io_c_24, pin_io_c_23, pin_io_c_22, pin_io_c_18, pin_io_c_14, 
        pin_io_c_13, pin_io_c_12, C_8_c;
    wire [15:0]spi_cmd_r;   // c:/s_links/sources/mcm_top.v(74[27:36])
    wire [7:0]spi_addr_r;   // c:/s_links/sources/mcm_top.v(75[28:38])
    wire [39:0]spi_data_r;   // c:/s_links/sources/mcm_top.v(76[22:32])
    
    wire spi_data_valid_r;
    wire [15:0]spi_cmd;   // c:/s_links/sources/mcm_top.v(79[27:34])
    wire [39:0]spi_data_out_r;   // c:/s_links/sources/mcm_top.v(81[22:36])
    wire [13:0]cs_decoded;   // c:/s_links/sources/mcm_top.v(84[43:53])
    
    wire n4;
    wire [6:0]quad_a;   // c:/s_links/sources/mcm_top.v(89[31:37])
    wire [6:0]quad_b;   // c:/s_links/sources/mcm_top.v(90[31:37])
    wire [6:0]pwm_out;   // c:/s_links/sources/mcm_top.v(96[31:38])
    wire [3:0]uart_slot_en;   // c:/s_links/sources/mcm_top.v(99[37:49])
    
    wire EM_STOP, VCC_net, spi_cmd_valid, spi_addr_valid, spi_data_valid, 
        clk_100k_enable_1, n26521, n29977, n29575, n12435, n23409, 
        n23722, n9;
    wire [13:0]cs_decoded_13__N_752;
    wire [12:0]status_cntr;   // c:/s_links/sources/status_led.v(37[32:43])
    
    wire pwm, n26243, pwm_N_898, clk_enable_263, clk_enable_638, n7164, 
        pwm_N_896, n2, n5, n29994, n4_adj_7388, n16, n23555;
    wire [39:0]spi_data_out_r_39__N_770;
    
    wire spi_data_out_r_39__N_810;
    wire [1:0]quad_homing;   // c:/s_links/sources/quad_decoder.v(40[19:30])
    wire [31:0]quad_count;   // c:/s_links/sources/quad_decoder.v(43[29:39])
    wire [31:0]quad_buffer;   // c:/s_links/sources/quad_decoder.v(44[29:40])
    
    wire quad_set_valid_N_1158, n11008;
    wire [39:0]spi_data_out_r_39__N_1083;
    wire [39:0]spi_data_out_r_39__N_934;
    
    wire spi_data_out_r_39__N_1163, spi_data_out_r_39__N_974, clk_enable_161, 
        n1, clk_enable_761, n29991, n29998, n30220, n7163, n23978, 
        n26207;
    wire [1:0]quad_homing_adj_7777;   // c:/s_links/sources/quad_decoder.v(40[19:30])
    
    wire quad_set_valid_N_1393, n18, n24700, n28524, n30110;
    wire [39:0]spi_data_out_r_39__N_1169;
    
    wire spi_data_out_r_39__N_1398, spi_data_out_r_39__N_1209, n23248, 
        n23610;
    wire [1:0]quad_homing_adj_7815;   // c:/s_links/sources/quad_decoder.v(40[19:30])
    wire [31:0]quad_count_adj_7816;   // c:/s_links/sources/quad_decoder.v(43[29:39])
    wire [31:0]quad_buffer_adj_7817;   // c:/s_links/sources/quad_decoder.v(44[29:40])
    wire [39:0]spi_data_out_r_39__N_1553;
    wire [39:0]spi_data_out_r_39__N_1404;
    
    wire spi_data_out_r_39__N_1633, spi_data_out_r_39__N_1444, n29997, 
        n29993, n28, n29996, clk_enable_38;
    wire [1:0]quad_homing_adj_7853;   // c:/s_links/sources/quad_decoder.v(40[19:30])
    
    wire n6747, n22554;
    wire [39:0]spi_data_out_r_39__N_1639;
    
    wire spi_data_out_r_39__N_1868, spi_data_out_r_39__N_1679, n1_adj_7459, 
        n6649, n18_adj_7460, n16_adj_7461, n5_adj_7462, n3;
    wire [1:0]quad_homing_adj_7891;   // c:/s_links/sources/quad_decoder.v(40[19:30])
    wire [31:0]quad_count_adj_7892;   // c:/s_links/sources/quad_decoder.v(43[29:39])
    wire [31:0]quad_buffer_adj_7893;   // c:/s_links/sources/quad_decoder.v(44[29:40])
    
    wire n23732, quad_set_valid_N_2098, n27095, n26497;
    wire [39:0]spi_data_out_r_39__N_2023;
    wire [39:0]spi_data_out_r_39__N_1874;
    
    wire spi_data_out_r_39__N_2103, spi_data_out_r_39__N_1914, n26119;
    wire [1:0]quad_homing_adj_7929;   // c:/s_links/sources/quad_decoder.v(40[19:30])
    wire [31:0]quad_count_adj_7930;   // c:/s_links/sources/quad_decoder.v(43[29:39])
    wire [31:0]quad_buffer_adj_7931;   // c:/s_links/sources/quad_decoder.v(44[29:40])
    
    wire quad_set_valid_N_2333, n26113;
    wire [39:0]spi_data_out_r_39__N_2258;
    wire [39:0]spi_data_out_r_39__N_2109;
    
    wire spi_data_out_r_39__N_2338, spi_data_out_r_39__N_2149, n19, n26107, 
        n18440, clk_enable_259;
    wire [1:0]quad_homing_adj_7967;   // c:/s_links/sources/quad_decoder.v(40[19:30])
    wire [31:0]quad_count_adj_7968;   // c:/s_links/sources/quad_decoder.v(43[29:39])
    wire [31:0]quad_buffer_adj_7969;   // c:/s_links/sources/quad_decoder.v(44[29:40])
    
    wire n26091, n26089, n23537;
    wire [39:0]spi_data_out_r_39__N_2493;
    wire [39:0]spi_data_out_r_39__N_2344;
    
    wire spi_data_out_r_39__N_2573, spi_data_out_r_39__N_2384, n22, n24169, 
        n21, clk_enable_23, clk_enable_759, n6651, n23916, n20647, 
        clear_intrpt;
    wire [39:0]spi_data_out_r_39__N_2579;
    
    wire intrpt_out_N_2642, clear_intrpt_adj_7661, n27015, clear_intrpt_N_2717;
    wire [39:0]spi_data_out_r_39__N_2650;
    
    wire n27013, intrpt_out_N_2713, clear_intrpt_adj_7662, clk_enable_227, 
        n2109, clear_intrpt_N_2788;
    wire [39:0]spi_data_out_r_39__N_2721;
    
    wire intrpt_out_N_2784, clear_intrpt_adj_7663, clear_intrpt_N_2859;
    wire [39:0]spi_data_out_r_39__N_2792;
    
    wire intrpt_out_N_2855, clear_intrpt_adj_7664, clear_intrpt_N_2930;
    wire [39:0]spi_data_out_r_39__N_2863;
    
    wire intrpt_out_N_2926, clear_intrpt_adj_7665, clear_intrpt_N_3001;
    wire [39:0]spi_data_out_r_39__N_2934;
    
    wire intrpt_out_N_2997, clear_intrpt_adj_7666, n57, clear_intrpt_N_3072;
    wire [39:0]spi_data_out_r_39__N_3005;
    
    wire intrpt_out_N_3068, pwm_out_N_3169, pwm_out_N_3153, n1_adj_7667, 
        n1_adj_7668, n1_adj_7669;
    wire [2:0]n31089;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    wire reset_r, digital_output_r, NSL, n47, n21_adj_7670, n26957, 
        n13, reset_r_N_4129, n6590, n26947;
    wire [39:0]spi_data_out_r_39__N_3825;
    
    wire spi_data_out_r_39__N_3865, reset_r_adj_7671, digital_output_r_adj_7672, 
        NSL_adj_7673;
    wire [51:0]SLO_buf_adj_8127;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire ENC_O_N_4469, OW_ID_N_4461, OW_ID_N_4467, n9_adj_7674, n28260;
    wire [39:0]spi_data_out_r_39__N_4419;
    wire [39:0]spi_data_out_r_39__N_4168;
    
    wire spi_data_out_r_39__N_4505, spi_data_out_r_39__N_4208, n2193, 
        n14;
    wire [2:0]n31091;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    wire reset_r_adj_7676, digital_output_r_adj_7677, NSL_adj_7678, ENC_O_N_4812, 
        OW_ID_N_4804, OW_ID_N_4810, n26873;
    wire [39:0]spi_data_out_r_39__N_4511;
    
    wire spi_data_out_r_39__N_4848, spi_data_out_r_39__N_4551, reset_r_adj_7679, 
        digital_output_r_adj_7680, NSL_adj_7681, n25979;
    wire [51:0]SLO_buf_adj_8193;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire ENC_O_N_5155, OW_ID_N_5147, OW_ID_N_5153, n1_adj_7712, n29995;
    wire [39:0]spi_data_out_r_39__N_5105;
    wire [39:0]spi_data_out_r_39__N_4854;
    
    wire spi_data_out_r_39__N_5191, spi_data_out_r_39__N_4894, reset_r_adj_7713, 
        digital_output_r_adj_7714, NSL_adj_7715, ENC_O_N_5498, OW_ID_N_5490, 
        OW_ID_N_5496, n26821, n28384, n26819, n25943, n25941, n30007, 
        n47_adj_7716;
    wire [39:0]spi_data_out_r_39__N_5197;
    
    wire spi_data_out_r_39__N_5534, spi_data_out_r_39__N_5237, reset_r_adj_7717, 
        digital_output_r_adj_7718, NSL_adj_7719, ENC_O_N_5841, OW_ID_N_5833, 
        OW_ID_N_5839, n30102, n26435, n25923, n26779;
    wire [39:0]spi_data_out_r_39__N_5540;
    
    wire spi_data_out_r_39__N_5877, spi_data_out_r_39__N_5580, reset_r_adj_7720, 
        digital_output_r_adj_7721, NSL_adj_7722, ENC_O_N_6184, OW_ID_N_6176, 
        OW_ID_N_6182, n25893, n25889, n25885, n25881, n25877, n25873, 
        n25869, n23148, clk_enable_254, n28486, n25859, n18654;
    wire [39:0]spi_data_out_r_39__N_5883;
    
    wire spi_data_out_r_39__N_6220, spi_data_out_r_39__N_5923, n1_adj_7723, 
        mode, Phase_r, mode_adj_7724, pwm_out_1, pwm_out_1_N_6306, 
        clk_enable_898, clk_enable_639, clk_enable_315, mode_adj_7725, 
        Phase_1_r, Phase_2_r, Phase_3_r, Phase_4_r;
    wire [11:0]pwm_duty_1_adj_8329;   // c:/s_links/sources/slot_cards/shutter_4.v(55[38:48])
    wire [11:0]pwm_duty_2_adj_8330;   // c:/s_links/sources/slot_cards/shutter_4.v(56[38:48])
    wire [11:0]pwm_duty_3_adj_8331;   // c:/s_links/sources/slot_cards/shutter_4.v(57[38:48])
    
    wire clk_enable_641, n28328, n5_adj_7726, pwm_out_1_N_6491, pwm_out_2_N_6511, 
        pwm_out_3_N_6530, pwm_out_4_N_6549, clk_enable_388, clk_enable_683, 
        clk_enable_684, clk_enable_727, clk_enable_687, mode_adj_7727, 
        TX_IN_N_6565, mode_adj_7728, mode_adj_7729, tx_N_6586, spi_mosi_oe, 
        spi_mosi_o, spi_miso_oe, spi_miso_o, spi_clk_oe, spi_clk_o, 
        spi_mosi_i, spi_miso_i, clk_enable_256, n47_adj_7730, n30098, 
        clk_enable_627, n25801, clk_enable_32, clk_enable_260, clk_enable_255, 
        clk_enable_253, clk_enable_245, clk_enable_244, clk_enable_749, 
        clk_enable_738, clk_enable_226, clk_enable_652, clk_enable_235, 
        clk_enable_232, clk_enable_234, clk_enable_15, n30095, n30094, 
        n28358, clk_enable_211, clk_enable_488, clk_enable_842, clk_enable_520, 
        clk_enable_807, clk_enable_180, clk_enable_22, n10696, n30091, 
        n30090, clk_enable_757, clk_enable_320, clk_enable_595, n47_adj_7731, 
        n29976, n29967, n8, n7, n25741, n47_adj_7732, n30087, 
        n25739, n26633, n25358, n26621, n29944, n29943, n25721, 
        n30083, n30004, n30082, n30080, n25699, n28544, n28476, 
        n30219, n25347, n30075, clk_enable_12, n29481, n26569, n24593, 
        n25643, clk_enable_222, n25212, n4_adj_7733, n30071, n30070, 
        n26545, n23526, n24066, n28402, n25223, n29992, n32, n47_adj_7734, 
        clk_enable_28, n29990, n30064, n30062, n25571, n26327, n30058, 
        n25547, n23609, n30055, clk_enable_242, n47_adj_7735, clk_enable_695, 
        n12467, n28340, n28562, n28561, n28560, n28559, n28558, 
        clk_enable_959, n30052, n30050, n7166, n7167, n7170, n11608, 
        n7177, n11013, n28557, n11609, n10500, n28556, n7198, 
        n7201, pin_io_out_69, pin_io_out_65, pin_io_out_59, pin_io_out_55, 
        pin_io_out_49, pin_io_out_45, pin_io_out_40, pin_io_out_39, 
        pin_io_out_35, pin_io_out_29, pin_io_out_25, pin_io_out_19, 
        pin_io_out_15, pin_io_out_9, pin_io_out_8, pin_io_out_6, pin_io_out_5, 
        pin_io_out_4, pin_io_out_3, pin_io_out_2, pin_io_out_1, n7258, 
        n7262, n7266, n7269, n7273, n7277, n28555, n30049, n28554, 
        clk_enable_1105, n30047, clk_enable_613, n11606, n28553, n28552, 
        n28551, n30235, n28550, n28549, n29999, n28548, clk_enable_1107, 
        n28547, n24588, n28546, n6, n30045, n30044, n30214, n30213, 
        n30210, n19_adj_7736, n20, n21_adj_7737, n30043, n30209, 
        n30203, n30199, n30198, n30188, n30185, n30041, n30039, 
        n30035, n30180, n30175, n31069, n30031, n30165, n30028, 
        n30027, n30023, n30155, n30218, n30151, n30149, n30020, 
        n30019, n30146, n30144, n30143, n30138, n30134, n30129, 
        n30018, n30125, n30122, clk_enable_686, clk_enable_178, n29594, 
        n30120, n30118, n30013;
    
    VHI i2 (.Z(VCC_net));
    OSCH OSCH_inst (.STDBY(GND_net), .OSC(clk)) /* synthesis syn_instantiated=1 */ ;
    defparam OSCH_inst.NOM_FREQ = "38.00";
    BB BBspi_mosi (.I(spi_mosi_o), .T(spi_mosi_oe), .B(spi_mosi), .O(spi_mosi_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=15, LSE_LLINE=162, LSE_RLINE=176 */ ;   // c:/s_links/sources/config_hex/ip/spi_slave_efb.v(39[8:82])
    BB BBspi_miso (.I(spi_miso_o), .T(spi_miso_oe), .B(spi_miso), .O(spi_miso_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=15, LSE_LLINE=162, LSE_RLINE=176 */ ;   // c:/s_links/sources/config_hex/ip/spi_slave_efb.v(41[8:82])
    BB BBspi_clk (.I(spi_clk_o), .T(spi_clk_oe), .B(spi_clk), .O(spi_clk_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=15, LSE_LLINE=162, LSE_RLINE=176 */ ;   // c:/s_links/sources/config_hex/ip/spi_slave_efb.v(43[8:77])
    \shutter(UART_ADDRESS_WIDTH=4)  \shutter_ins_0..u_shutter  (.clk(clk), 
            .clk_enable_22(clk_enable_22), .n6590(n6590), .Phase_4_r(Phase_4_r), 
            .clk_enable_244(clk_enable_244), .n30185(n30185), .n28546(n28546), 
            .\spi_cmd_r[3] (spi_cmd_r[3]), .n30064(n30064), .n23916(n23916), 
            .n26435(n26435), .clk_enable_695(clk_enable_695), .pwm_duty_2({pwm_duty_2_adj_8330}), 
            .clk_enable_226(clk_enable_226), .\spi_data_r[0] (spi_data_r[0]), 
            .n29998(n29998), .pwm_duty_1({pwm_duty_1_adj_8329}), .clk_enable_652(clk_enable_652), 
            .pwm_duty_3({pwm_duty_3_adj_8331}), .clk_enable_738(clk_enable_738), 
            .clk_enable_749(clk_enable_749), .\spi_data_r[11] (spi_data_r[11]), 
            .\spi_data_r[10] (spi_data_r[10]), .\spi_data_r[9] (spi_data_r[9]), 
            .\spi_data_r[8] (spi_data_r[8]), .\spi_data_r[7] (spi_data_r[7]), 
            .\spi_data_r[6] (spi_data_r[6]), .\spi_data_r[5] (spi_data_r[5]), 
            .Phase_1_r(Phase_1_r), .n28548(n28548), .\spi_data_r[4] (spi_data_r[4]), 
            .\spi_data_r[3] (spi_data_r[3]), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[1] (spi_data_r[1]), .GND_net(GND_net), .Phase_2_r(Phase_2_r), 
            .n28552(n28552), .Phase_3_r(Phase_3_r), .n28553(n28553), .mode(mode_adj_7725), 
            .clk_enable_245(clk_enable_245), .clk_enable_613(clk_enable_613), 
            .n6747(n6747), .\spi_cmd_r[2] (spi_cmd_r[2]), .\spi_cmd_r[0] (spi_cmd_r[0]), 
            .\spi_addr_r[2] (spi_addr_r[2]), .\spi_addr_r[6] (spi_addr_r[6]), 
            .n26243(n26243), .\spi_data_r[17] (spi_data_r[17]), .\spi_data_r[16] (spi_data_r[16]), 
            .n26521(n26521), .n21(n21_adj_7737), .n19(n19_adj_7736), .n20(n20), 
            .n26545(n26545), .\spi_addr_r[4] (spi_addr_r[4]), .n26497(n26497), 
            .n26569(n26569), .pwm_out_4_N_6549(pwm_out_4_N_6549), .pwm_out_1_N_6491(pwm_out_1_N_6491), 
            .pwm_out_3_N_6530(pwm_out_3_N_6530), .NSL(NSL), .n30058(n30058), 
            .n25347(n25347), .\pwm_out[0] (pwm_out[0]), .mode_adj_660(mode), 
            .pwm_out_1(pwm_out_1), .mode_adj_661(mode_adj_7724), .reset_r(reset_r), 
            .n30043(n30043), .n25223(n25223), .n4(n4_adj_7733), .mode_adj_662({n31089}), 
            .digital_output_r(digital_output_r), .n23148(n23148), .Phase_r(Phase_r), 
            .n24593(n24593), .UC_TXD0_c(UC_TXD0_c), .n23409(n23409), .\uart_slot_en[3] (uart_slot_en[3]), 
            .n30125(n30125), .\cs_decoded[0] (cs_decoded[0]), .n11013(n11013), 
            .n30018(n30018), .n8(n8), .n23722(n23722), .n23555(n23555), 
            .n30129(n30129), .n30052(n30052), .n24588(n24588), .pwm_out_2_N_6511(pwm_out_2_N_6511), 
            .n23610(n23610), .clk_enable_1105(clk_enable_1105), .n6651(n6651), 
            .clk_enable_1107(clk_enable_1107), .n6649(n6649), .n10500(n10500), 
            .n7198(n7198), .n7177(n7177), .n7201(n7201), .n30134(n30134), 
            .n11609(n11609), .n30175(n30175), .n11606(n11606), .n11608(n11608), 
            .n11008(n11008)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(498[3] 530[2])
    IB C_8_pad (.I(C_8), .O(C_8_c));   // c:/s_links/sources/mcm_top.v(46[24:27])
    IB pin_io_pad_12 (.I(pin_io[12]), .O(pin_io_c_12));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_13 (.I(pin_io[13]), .O(pin_io_c_13));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_14 (.I(pin_io[14]), .O(pin_io_c_14));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_18 (.I(pin_io[18]), .O(pin_io_c_18));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_22 (.I(pin_io[22]), .O(pin_io_c_22));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_23 (.I(pin_io[23]), .O(pin_io_c_23));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_24 (.I(pin_io[24]), .O(pin_io_c_24));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_28 (.I(pin_io[28]), .O(pin_io_c_28));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_32 (.I(pin_io[32]), .O(pin_io_c_32));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_33 (.I(pin_io[33]), .O(pin_io_c_33));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_34 (.I(pin_io[34]), .O(pin_io_c_34));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_38 (.I(pin_io[38]), .O(pin_io_c_38));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_42 (.I(pin_io[42]), .O(pin_io_c_42));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_43 (.I(pin_io[43]), .O(pin_io_c_43));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_44 (.I(pin_io[44]), .O(pin_io_c_44));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_48 (.I(pin_io[48]), .O(pin_io_c_48));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_52 (.I(pin_io[52]), .O(pin_io_c_52));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_53 (.I(pin_io[53]), .O(pin_io_c_53));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_54 (.I(pin_io[54]), .O(pin_io_c_54));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_58 (.I(pin_io[58]), .O(pin_io_c_58));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_62 (.I(pin_io[62]), .O(pin_io_c_62));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_63 (.I(pin_io[63]), .O(pin_io_c_63));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_64 (.I(pin_io[64]), .O(pin_io_c_64));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB pin_io_pad_68 (.I(pin_io[68]), .O(pin_io_c_68));   // c:/s_links/sources/mcm_top.v(36[51:57])
    IB UC_TXD0_pad (.I(UC_TXD0), .O(UC_TXD0_c));   // c:/s_links/sources/mcm_top.v(32[27:34])
    IB spi_scsn_pad (.I(spi_scsn), .O(spi_scsn_c));   // c:/s_links/sources/mcm_top.v(29[27:35])
    IB CS_READY_pad (.I(CS_READY), .O(CS_READY_c));   // c:/s_links/sources/mcm_top.v(23[24:32])
    IB cs_pad_0 (.I(cs[0]), .O(cs_c_0));   // c:/s_links/sources/mcm_top.v(19[37:39])
    IB cs_pad_1 (.I(cs[1]), .O(cs_c_1));   // c:/s_links/sources/mcm_top.v(19[37:39])
    IB cs_pad_2 (.I(cs[2]), .O(cs_c_2));   // c:/s_links/sources/mcm_top.v(19[37:39])
    IB cs_pad_3 (.I(cs[3]), .O(cs_c_3));   // c:/s_links/sources/mcm_top.v(19[37:39])
    IB cs_pad_4 (.I(cs[4]), .O(cs_c_4));   // c:/s_links/sources/mcm_top.v(19[37:39])
    IB resetn_pad (.I(resetn), .O(resetn_c));   // c:/s_links/sources/mcm_top.v(17[27:33])
    IB clk_in_pad (.I(clk_in), .O(clk_in_c));   // c:/s_links/sources/mcm_top.v(16[27:33])
    OBZ C_7_pad (.I(UC_TXD0_c), .T(tx_N_6586), .O(C_7));   // c:/s_links/sources/slot_cards/peizo_elliptec.v(30[8:10])
    OBZ pin_io_pad_0 (.I(n23610), .T(n23609), .O(pin_io[0]));
    OBZ pin_io_pad_7 (.I(n25347), .T(n23609), .O(pin_io[7]));
    OBZ pin_io_pad_10 (.I(VCC_net), .T(n30041), .O(pin_io[10]));   // c:/s_links/sources/slot_cards/stepper.v(70[8:10])
    OBZ pin_io_pad_11 (.I(reset_r_adj_7671), .T(n7277), .O(pin_io[11]));   // c:/s_links/sources/slot_cards/stepper.v(71[8:13])
    OBZ pin_io_pad_16 (.I(cs_decoded[2]), .T(n7277), .O(pin_io[16]));   // c:/s_links/sources/slot_cards/stepper.v(75[8:14])
    OBZ pin_io_pad_17 (.I(NSL_adj_7673), .T(n30041), .O(pin_io[17]));   // c:/s_links/sources/slot_cards/stepper.v(76[8:15])
    OBZ pin_io_pad_20 (.I(VCC_net), .T(n5_adj_7726), .O(pin_io[20]));   // c:/s_links/sources/slot_cards/stepper.v(70[8:10])
    OBZ pin_io_pad_21 (.I(reset_r_adj_7676), .T(n7273), .O(pin_io[21]));   // c:/s_links/sources/slot_cards/stepper.v(71[8:13])
    OBZ pin_io_pad_26 (.I(cs_decoded[4]), .T(n7273), .O(pin_io[26]));   // c:/s_links/sources/slot_cards/stepper.v(75[8:14])
    OBZ pin_io_pad_27 (.I(NSL_adj_7678), .T(n5_adj_7726), .O(pin_io[27]));   // c:/s_links/sources/slot_cards/stepper.v(76[8:15])
    OBZ pin_io_pad_30 (.I(n7170), .T(n7166), .O(pin_io[30]));
    OBZ pin_io_pad_31 (.I(reset_r_adj_7679), .T(n7269), .O(pin_io[31]));   // c:/s_links/sources/slot_cards/stepper.v(71[8:13])
    OBZ pin_io_pad_36 (.I(cs_decoded[6]), .T(n7269), .O(pin_io[36]));   // c:/s_links/sources/slot_cards/stepper.v(75[8:14])
    OBZ pin_io_pad_37 (.I(n7167), .T(n7166), .O(pin_io[37]));
    OBZ pin_io_pad_41 (.I(reset_r_adj_7713), .T(n7266), .O(pin_io[41]));   // c:/s_links/sources/slot_cards/stepper.v(71[8:13])
    OBZ pin_io_pad_46 (.I(cs_decoded[8]), .T(n7266), .O(pin_io[46]));   // c:/s_links/sources/slot_cards/stepper.v(75[8:14])
    OBZ pin_io_pad_47 (.I(NSL_adj_7715), .T(n30180), .O(pin_io[47]));   // c:/s_links/sources/slot_cards/stepper.v(76[8:15])
    OBZ pin_io_pad_50 (.I(VCC_net), .T(n30047), .O(pin_io[50]));   // c:/s_links/sources/slot_cards/stepper.v(70[8:10])
    OBZ pin_io_pad_51 (.I(reset_r_adj_7717), .T(n7262), .O(pin_io[51]));   // c:/s_links/sources/slot_cards/stepper.v(71[8:13])
    OBZ pin_io_pad_56 (.I(cs_decoded[10]), .T(n7262), .O(pin_io[56]));   // c:/s_links/sources/slot_cards/stepper.v(75[8:14])
    OBZ pin_io_pad_57 (.I(NSL_adj_7719), .T(n30047), .O(pin_io[57]));   // c:/s_links/sources/slot_cards/stepper.v(76[8:15])
    OBZ pin_io_pad_60 (.I(VCC_net), .T(n30165), .O(pin_io[60]));   // c:/s_links/sources/slot_cards/stepper.v(70[8:10])
    OBZ pin_io_pad_61 (.I(reset_r_adj_7720), .T(n7258), .O(pin_io[61]));   // c:/s_links/sources/slot_cards/stepper.v(71[8:13])
    OBZ pin_io_pad_66 (.I(cs_decoded[12]), .T(n7258), .O(pin_io[66]));   // c:/s_links/sources/slot_cards/stepper.v(75[8:14])
    OBZ pin_io_pad_67 (.I(NSL_adj_7722), .T(n30165), .O(pin_io[67]));   // c:/s_links/sources/slot_cards/stepper.v(76[8:15])
    OBZ UC_RXD0_pad (.I(n23248), .T(n25358), .O(UC_RXD0));
    OB MAX3421_CS_pad (.I(MAX3421_CS_c), .O(MAX3421_CS));   // c:/s_links/sources/mcm_top.v(22[24:34])
    OB FLASH_CS_pad (.I(FLASH_CS_c), .O(FLASH_CS));   // c:/s_links/sources/mcm_top.v(21[24:32])
    OB intrpt_out_pad_0 (.I(intrpt_out_c_0), .O(intrpt_out[0]));   // c:/s_links/sources/mcm_top.v(20[36:46])
    OB intrpt_out_pad_1 (.I(intrpt_out_c_1), .O(intrpt_out[1]));   // c:/s_links/sources/mcm_top.v(20[36:46])
    OB intrpt_out_pad_2 (.I(intrpt_out_c_2), .O(intrpt_out[2]));   // c:/s_links/sources/mcm_top.v(20[36:46])
    OB intrpt_out_pad_3 (.I(intrpt_out_c_3), .O(intrpt_out[3]));   // c:/s_links/sources/mcm_top.v(20[36:46])
    OB intrpt_out_pad_4 (.I(intrpt_out_c_4), .O(intrpt_out[4]));   // c:/s_links/sources/mcm_top.v(20[36:46])
    OB intrpt_out_pad_5 (.I(intrpt_out_c_5), .O(intrpt_out[5]));   // c:/s_links/sources/mcm_top.v(20[36:46])
    OB intrpt_out_pad_6 (.I(intrpt_out_c_6), .O(intrpt_out[6]));   // c:/s_links/sources/mcm_top.v(20[36:46])
    OB led_sw_pad (.I(led_sw_c), .O(led_sw));   // c:/s_links/sources/mcm_top.v(18[24:30])
    BB pin_io_pad_1 (.I(n25223), .T(n11609), .B(pin_io[1]), .O(pin_io_out_1));
    BB pin_io_pad_2 (.I(n7201), .T(n30125), .B(pin_io[2]), .O(pin_io_out_2));
    BB pin_io_pad_3 (.I(n7198), .T(n30125), .B(pin_io[3]), .O(pin_io_out_3));
    BB pin_io_pad_4 (.I(n10500), .T(n11608), .B(pin_io[4]), .O(pin_io_out_4));
    BB pin_io_pad_5 (.I(n23148), .T(n24593), .B(pin_io[5]), .O(pin_io_out_5));
    BB pin_io_pad_6 (.I(n11013), .T(n23555), .B(pin_io[6]), .O(pin_io_out_6));
    BB pin_io_pad_8 (.I(n7177), .T(n30125), .B(pin_io[8]), .O(pin_io_out_8));
    BB pin_io_pad_9 (.I(n24588), .T(n11606), .B(pin_io[9]), .O(pin_io_out_9));
    BB pin_io_pad_15 (.I(OW_ID_N_4461), .T(OW_ID_N_4467), .B(pin_io[15]), 
       .O(pin_io_out_15));   // c:/s_links/sources/slot_cards/stepper.v(90[8:13])
    BB pin_io_pad_19 (.I(n30098), .T(ENC_O_N_4469), .B(pin_io[19]), .O(pin_io_out_19));   // c:/s_links/sources/slot_cards/stepper.v(80[8:13])
    BB pin_io_pad_25 (.I(OW_ID_N_4804), .T(OW_ID_N_4810), .B(pin_io[25]), 
       .O(pin_io_out_25));   // c:/s_links/sources/slot_cards/stepper.v(90[8:13])
    BB pin_io_pad_29 (.I(n30110), .T(ENC_O_N_4812), .B(pin_io[29]), .O(pin_io_out_29));   // c:/s_links/sources/slot_cards/stepper.v(80[8:13])
    BB pin_io_pad_35 (.I(OW_ID_N_5147), .T(OW_ID_N_5153), .B(pin_io[35]), 
       .O(pin_io_out_35));   // c:/s_links/sources/slot_cards/stepper.v(90[8:13])
    BB pin_io_pad_39 (.I(n30188), .T(ENC_O_N_5155), .B(pin_io[39]), .O(pin_io_out_39));   // c:/s_links/sources/slot_cards/stepper.v(80[8:13])
    BB pin_io_pad_40 (.I(n7164), .T(n7163), .B(pin_io[40]), .O(pin_io_out_40));
    BB pin_io_pad_45 (.I(OW_ID_N_5490), .T(OW_ID_N_5496), .B(pin_io[45]), 
       .O(pin_io_out_45));   // c:/s_links/sources/slot_cards/stepper.v(90[8:13])
    BB pin_io_pad_49 (.I(n30146), .T(ENC_O_N_5498), .B(pin_io[49]), .O(pin_io_out_49));   // c:/s_links/sources/slot_cards/stepper.v(80[8:13])
    BB pin_io_pad_55 (.I(OW_ID_N_5833), .T(OW_ID_N_5839), .B(pin_io[55]), 
       .O(pin_io_out_55));   // c:/s_links/sources/slot_cards/stepper.v(90[8:13])
    BB pin_io_pad_59 (.I(n30149), .T(ENC_O_N_5841), .B(pin_io[59]), .O(pin_io_out_59));   // c:/s_links/sources/slot_cards/stepper.v(80[8:13])
    BB pin_io_pad_65 (.I(OW_ID_N_6176), .T(OW_ID_N_6182), .B(pin_io[65]), 
       .O(pin_io_out_65));   // c:/s_links/sources/slot_cards/stepper.v(90[8:13])
    BB pin_io_pad_69 (.I(n30143), .T(ENC_O_N_6184), .B(pin_io[69]), .O(pin_io_out_69));   // c:/s_links/sources/slot_cards/stepper.v(80[8:13])
    LUT4 i1847_4_lut (.A(spi_addr_valid), .B(n30080), .C(spi_cmd_valid), 
         .D(spi_data_valid), .Z(clk_enable_161)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;
    defparam i1847_4_lut.init = 16'hcdcc;
    LUT4 i23844_4_lut (.A(Phase_4_r), .B(spi_data_r[0]), .C(spi_data_r[1]), 
         .D(spi_data_r[2]), .Z(n28546)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i23844_4_lut.init = 16'hcaaa;
    VLO i1 (.Z(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i23845_4_lut (.A(digital_output_r), .B(spi_data_r[0]), .C(n25571), 
         .D(n23916), .Z(n28547)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i23845_4_lut.init = 16'hcaaa;
    \intrpt_ctrl(DEV_ID=1)  \intrpt_ins_1..u_intrpt_ctrl  (.clear_intrpt(clear_intrpt_adj_7661), 
            .clk(clk), .n30185(n30185), .clear_intrpt_N_2717(clear_intrpt_N_2717), 
            .\spi_data_out_r_39__N_2650[0] (spi_data_out_r_39__N_2650[0]), 
            .\pin_intrpt[3] (pin_intrpt[3]), .\pin_intrpt[5] (pin_intrpt[5]), 
            .\pin_intrpt[4] (pin_intrpt[4]), .intrpt_out_c_1(intrpt_out_c_1), 
            .intrpt_out_N_2713(intrpt_out_N_2713), .n31069(n31069), .\spi_data_out_r_39__N_2650[2] (spi_data_out_r_39__N_2650[2]), 
            .\spi_data_out_r_39__N_2650[1] (spi_data_out_r_39__N_2650[1])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(294[3] 315[2])
    \intrpt_ctrl(DEV_ID=2)  \intrpt_ins_2..u_intrpt_ctrl  (.clk(clk), .n30185(n30185), 
            .\spi_data_out_r_39__N_2721[0] (spi_data_out_r_39__N_2721[0]), 
            .\pin_intrpt[6] (pin_intrpt[6]), .clear_intrpt(clear_intrpt_adj_7662), 
            .clear_intrpt_N_2788(clear_intrpt_N_2788), .\pin_intrpt[8] (pin_intrpt[8]), 
            .\pin_intrpt[7] (pin_intrpt[7]), .intrpt_out_c_2(intrpt_out_c_2), 
            .intrpt_out_N_2784(intrpt_out_N_2784), .n31069(n31069), .\spi_data_out_r_39__N_2721[2] (spi_data_out_r_39__N_2721[2]), 
            .\spi_data_out_r_39__N_2721[1] (spi_data_out_r_39__N_2721[1])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(294[3] 315[2])
    LUT4 i23846_4_lut (.A(Phase_1_r), .B(spi_data_r[0]), .C(spi_data_r[1]), 
         .D(spi_data_r[2]), .Z(n28548)) /* synthesis lut_function=(A (B+(C+(D)))+!A !((C+(D))+!B)) */ ;
    defparam i23846_4_lut.init = 16'haaac;
    LUT4 i23843_4_lut_then_4_lut (.A(cs_c_4), .B(cs_c_3), .C(cs_c_2), 
         .D(cs_c_0), .Z(n30219)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;
    defparam i23843_4_lut_then_4_lut.init = 16'h7fff;
    LUT4 i23847_4_lut (.A(digital_output_r_adj_7714), .B(spi_data_r[0]), 
         .C(n23916), .D(n25943), .Z(n28549)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i23847_4_lut.init = 16'hcaaa;
    LUT4 i23855_4_lut (.A(cs_decoded[12]), .B(cs_c_1), .C(n30235), .D(n30203), 
         .Z(n28557)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i23855_4_lut.init = 16'hfaca;
    LUT4 i23856_4_lut (.A(cs_decoded[10]), .B(cs_decoded_13__N_752[10]), 
         .C(cs_c_4), .D(n29977), .Z(n28558)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;
    defparam i23856_4_lut.init = 16'hccca;
    LUT4 i23857_4_lut (.A(cs_decoded[8]), .B(cs_decoded_13__N_752[10]), 
         .C(cs_c_4), .D(n29976), .Z(n28559)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;
    defparam i23857_4_lut.init = 16'hccca;
    LUT4 i23848_4_lut (.A(digital_output_r_adj_7721), .B(spi_data_r[0]), 
         .C(n23916), .D(n25923), .Z(n28550)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i23848_4_lut.init = 16'hcaaa;
    intrpt_ctrl \intrpt_ins_0..u_intrpt_ctrl  (.intrpt_out_c_0(intrpt_out_c_0), 
            .clk(clk), .intrpt_out_N_2642(intrpt_out_N_2642), .n31069(n31069), 
            .n30185(n30185), .\spi_data_out_r_39__N_2579[0] (spi_data_out_r_39__N_2579[0]), 
            .\pin_intrpt[0] (pin_intrpt[0]), .clear_intrpt(clear_intrpt), 
            .\spi_data_out_r_39__N_2579[2] (spi_data_out_r_39__N_2579[2]), 
            .\pin_intrpt[2] (pin_intrpt[2]), .\spi_data_out_r_39__N_2579[1] (spi_data_out_r_39__N_2579[1]), 
            .\pin_intrpt[1] (pin_intrpt[1]), .n30198(n30198), .n30019(n30019), 
            .n30013(n30013), .n30027(n30027)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(294[3] 315[2])
    LUT4 i23858_4_lut (.A(cs_decoded[6]), .B(cs_decoded_13__N_752[6]), .C(cs_c_4), 
         .D(n13), .Z(n28560)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;
    defparam i23858_4_lut.init = 16'hccca;
    LUT4 i23859_4_lut (.A(cs_decoded[4]), .B(cs_decoded_13__N_752[6]), .C(cs_c_4), 
         .D(n29967), .Z(n28561)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;
    defparam i23859_4_lut.init = 16'hccca;
    LUT4 i23860_4_lut (.A(pwm), .B(pwm_N_896), .C(pwm_N_898), .D(n12467), 
         .Z(n28562)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;
    defparam i23860_4_lut.init = 16'hccca;
    \intrpt_ctrl(DEV_ID=5)  \intrpt_ins_5..u_intrpt_ctrl  (.clear_intrpt(clear_intrpt_adj_7665), 
            .clk(clk), .n30185(n30185), .clear_intrpt_N_3001(clear_intrpt_N_3001), 
            .intrpt_out_c_5(intrpt_out_c_5), .intrpt_out_N_2997(intrpt_out_N_2997), 
            .n31069(n31069), .\spi_data_out_r_39__N_2934[0] (spi_data_out_r_39__N_2934[0]), 
            .\pin_intrpt[15] (pin_intrpt[15]), .\spi_data_out_r_39__N_2934[2] (spi_data_out_r_39__N_2934[2]), 
            .\pin_intrpt[17] (pin_intrpt[17]), .\spi_data_out_r_39__N_2934[1] (spi_data_out_r_39__N_2934[1]), 
            .\pin_intrpt[16] (pin_intrpt[16])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(294[3] 315[2])
    \intrpt_ctrl(DEV_ID=3)  \intrpt_ins_3..u_intrpt_ctrl  (.clk(clk), .n30185(n30185), 
            .\spi_data_out_r_39__N_2792[0] (spi_data_out_r_39__N_2792[0]), 
            .\pin_intrpt[9] (pin_intrpt[9]), .clear_intrpt(clear_intrpt_adj_7663), 
            .clear_intrpt_N_2859(clear_intrpt_N_2859), .\pin_intrpt[11] (pin_intrpt[11]), 
            .\pin_intrpt[10] (pin_intrpt[10]), .intrpt_out_c_3(intrpt_out_c_3), 
            .intrpt_out_N_2855(intrpt_out_N_2855), .n31069(n31069), .\spi_data_out_r_39__N_2792[2] (spi_data_out_r_39__N_2792[2]), 
            .\spi_data_out_r_39__N_2792[1] (spi_data_out_r_39__N_2792[1])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(294[3] 315[2])
    cs_decoder u_cs_decoder (.\cs_decoded[0] (cs_decoded[0]), .CS_READY_c(CS_READY_c), 
            .n28544(n28544), .FLASH_CS_c(FLASH_CS_c), .n30220(n30220), 
            .MAX3421_CS_c(MAX3421_CS_c), .cs_c_3(cs_c_3), .cs_c_2(cs_c_2), 
            .cs_c_4(cs_c_4), .cs_c_0(cs_c_0), .cs_c_1(cs_c_1), .n13(n13), 
            .\cs_decoded[12] (cs_decoded[12]), .n28557(n28557), .\cs_decoded[10] (cs_decoded[10]), 
            .n28558(n28558), .\cs_decoded[8] (cs_decoded[8]), .n28559(n28559), 
            .\cs_decoded[6] (cs_decoded[6]), .n28560(n28560), .\cs_decoded[4] (cs_decoded[4]), 
            .n28561(n28561), .n29575(n29575), .\cs_decoded_13__N_752[6] (cs_decoded_13__N_752[6]), 
            .\cs_decoded_13__N_752[0] (cs_decoded_13__N_752[0]), .n30203(n30203), 
            .\cs_decoded_13__N_752[10] (cs_decoded_13__N_752[10]), .n29967(n29967), 
            .\cs_decoded[2] (cs_decoded[2]), .n29976(n29976), .n29977(n29977), 
            .n30235(n30235)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(204[3] 212[2])
    LUT4 i23842_4_lut (.A(cs_decoded[0]), .B(cs_decoded_13__N_752[0]), .C(cs_c_4), 
         .D(n29575), .Z(n28544)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;
    defparam i23842_4_lut.init = 16'hccca;
    \quad_decoder(DEV_ID=1)  \quad_ins_1..u_quad_decoder  (.quad_homing({quad_homing_adj_7777}), 
            .clk(clk), .clk_enable_520(clk_enable_520), .n30185(n30185), 
            .\spi_data_r[0] (spi_data_r[0]), .\quad_a[1] (quad_a[1]), .\quad_b[1] (quad_b[1]), 
            .\spi_data_out_r_39__N_1169[0] (spi_data_out_r_39__N_1169[0]), 
            .\pin_intrpt[5] (pin_intrpt[5]), .GND_net(GND_net), .clk_enable_842(clk_enable_842), 
            .quad_set_valid_N_1393(quad_set_valid_N_1393), .spi_data_out_r_39__N_1209(spi_data_out_r_39__N_1209), 
            .spi_data_out_r_39__N_1398(spi_data_out_r_39__N_1398), .\spi_data_out_r_39__N_1169[31] (spi_data_out_r_39__N_1169[31]), 
            .\spi_data_out_r_39__N_1169[30] (spi_data_out_r_39__N_1169[30]), 
            .\spi_data_out_r_39__N_1169[29] (spi_data_out_r_39__N_1169[29]), 
            .\spi_data_out_r_39__N_1169[28] (spi_data_out_r_39__N_1169[28]), 
            .\spi_data_out_r_39__N_1169[27] (spi_data_out_r_39__N_1169[27]), 
            .\spi_data_out_r_39__N_1169[26] (spi_data_out_r_39__N_1169[26]), 
            .\spi_data_out_r_39__N_1169[25] (spi_data_out_r_39__N_1169[25]), 
            .\spi_data_out_r_39__N_1169[24] (spi_data_out_r_39__N_1169[24]), 
            .\spi_data_out_r_39__N_1169[23] (spi_data_out_r_39__N_1169[23]), 
            .\spi_data_out_r_39__N_1169[22] (spi_data_out_r_39__N_1169[22]), 
            .\spi_data_out_r_39__N_1169[21] (spi_data_out_r_39__N_1169[21]), 
            .\spi_data_out_r_39__N_1169[20] (spi_data_out_r_39__N_1169[20]), 
            .\spi_data_out_r_39__N_1169[19] (spi_data_out_r_39__N_1169[19]), 
            .\spi_data_out_r_39__N_1169[18] (spi_data_out_r_39__N_1169[18]), 
            .\spi_data_out_r_39__N_1169[17] (spi_data_out_r_39__N_1169[17]), 
            .\spi_data_out_r_39__N_1169[16] (spi_data_out_r_39__N_1169[16]), 
            .\spi_data_out_r_39__N_1169[15] (spi_data_out_r_39__N_1169[15]), 
            .\spi_data_out_r_39__N_1169[14] (spi_data_out_r_39__N_1169[14]), 
            .\spi_data_out_r_39__N_1169[13] (spi_data_out_r_39__N_1169[13]), 
            .\spi_data_out_r_39__N_1169[12] (spi_data_out_r_39__N_1169[12]), 
            .\spi_data_out_r_39__N_1169[11] (spi_data_out_r_39__N_1169[11]), 
            .\spi_data_out_r_39__N_1169[10] (spi_data_out_r_39__N_1169[10]), 
            .\spi_data_out_r_39__N_1169[9] (spi_data_out_r_39__N_1169[9]), 
            .\spi_data_out_r_39__N_1169[8] (spi_data_out_r_39__N_1169[8]), 
            .\spi_data_out_r_39__N_1169[7] (spi_data_out_r_39__N_1169[7]), 
            .\spi_data_out_r_39__N_1169[6] (spi_data_out_r_39__N_1169[6]), 
            .\spi_data_out_r_39__N_1169[5] (spi_data_out_r_39__N_1169[5]), 
            .\spi_data_out_r_39__N_1169[4] (spi_data_out_r_39__N_1169[4]), 
            .\spi_data_out_r_39__N_1169[3] (spi_data_out_r_39__N_1169[3]), 
            .\spi_data_out_r_39__N_1169[2] (spi_data_out_r_39__N_1169[2]), 
            .\spi_data_out_r_39__N_1169[1] (spi_data_out_r_39__N_1169[1]), 
            .\spi_data_r[1] (spi_data_r[1]), .n47(n47_adj_7735), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[3] (spi_data_r[3]), .\spi_data_r[4] (spi_data_r[4]), 
            .\spi_data_r[5] (spi_data_r[5]), .\spi_data_r[6] (spi_data_r[6]), 
            .\spi_data_r[7] (spi_data_r[7]), .\spi_data_r[8] (spi_data_r[8]), 
            .\spi_data_r[9] (spi_data_r[9]), .\spi_data_r[10] (spi_data_r[10]), 
            .\spi_data_r[11] (spi_data_r[11]), .\spi_data_r[12] (spi_data_r[12]), 
            .\spi_data_r[13] (spi_data_r[13]), .\spi_data_r[14] (spi_data_r[14]), 
            .\spi_data_r[15] (spi_data_r[15]), .\spi_data_r[16] (spi_data_r[16]), 
            .\spi_data_r[17] (spi_data_r[17]), .\spi_data_r[18] (spi_data_r[18]), 
            .\spi_data_r[19] (spi_data_r[19]), .\spi_data_r[20] (spi_data_r[20]), 
            .\spi_data_r[21] (spi_data_r[21]), .\spi_data_r[22] (spi_data_r[22]), 
            .\spi_data_r[23] (spi_data_r[23]), .\spi_data_r[24] (spi_data_r[24]), 
            .\spi_data_r[25] (spi_data_r[25]), .\spi_data_r[26] (spi_data_r[26]), 
            .\spi_data_r[27] (spi_data_r[27]), .\spi_data_r[28] (spi_data_r[28]), 
            .\spi_data_r[29] (spi_data_r[29]), .\spi_data_r[30] (spi_data_r[30]), 
            .\spi_data_r[31] (spi_data_r[31]), .n1(n1_adj_7668), .resetn_c(resetn_c)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(263[3] 283[2])
    LUT4 i23849_4_lut (.A(digital_output_r_adj_7718), .B(spi_data_r[0]), 
         .C(n27015), .D(n23916), .Z(n28551)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i23849_4_lut.init = 16'hcaaa;
    LUT4 i23850_4_lut (.A(Phase_2_r), .B(spi_data_r[0]), .C(spi_data_r[1]), 
         .D(spi_data_r[2]), .Z(n28552)) /* synthesis lut_function=(A (B+((D)+!C))+!A !(((D)+!C)+!B)) */ ;
    defparam i23850_4_lut.init = 16'haaca;
    LUT4 i23851_4_lut (.A(Phase_3_r), .B(spi_data_r[0]), .C(spi_data_r[1]), 
         .D(spi_data_r[2]), .Z(n28553)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !((C+!(D))+!B)) */ ;
    defparam i23851_4_lut.init = 16'hacaa;
    LUT4 i23852_4_lut (.A(digital_output_r_adj_7680), .B(spi_data_r[0]), 
         .C(n25859), .D(n28524), .Z(n28554)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;
    defparam i23852_4_lut.init = 16'hccac;
    LUT4 i23853_4_lut (.A(digital_output_r_adj_7672), .B(spi_data_r[0]), 
         .C(n25801), .D(n28524), .Z(n28555)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C))) */ ;
    defparam i23853_4_lut.init = 16'hccac;
    LUT4 i23854_4_lut (.A(digital_output_r_adj_7677), .B(spi_data_r[0]), 
         .C(n26119), .D(n23916), .Z(n28556)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;
    defparam i23854_4_lut.init = 16'hcacc;
    \quad_decoder(DEV_ID=6)  \quad_ins_6..u_quad_decoder  (.GND_net(GND_net), 
            .quad_count({quad_count_adj_7968}), .clk(clk), .n30185(n30185), 
            .\quad_a[6] (quad_a[6]), .\quad_b[6] (quad_b[6]), .\spi_data_out_r_39__N_2344[0] (spi_data_out_r_39__N_2344[0]), 
            .\spi_data_out_r_39__N_2493[0] (spi_data_out_r_39__N_2493[0]), 
            .quad_buffer({quad_buffer_adj_7969}), .\pin_intrpt[20] (pin_intrpt[20]), 
            .n30004(n30004), .spi_data_out_r_39__N_2384(spi_data_out_r_39__N_2384), 
            .spi_data_out_r_39__N_2573(spi_data_out_r_39__N_2573), .quad_homing({quad_homing_adj_7967}), 
            .clk_enable_639(clk_enable_639), .\spi_data_r[0] (spi_data_r[0]), 
            .clk_enable_898(clk_enable_898), .\spi_data_out_r_39__N_2344[31] (spi_data_out_r_39__N_2344[31]), 
            .\spi_data_out_r_39__N_2493[31] (spi_data_out_r_39__N_2493[31]), 
            .\spi_data_out_r_39__N_2344[30] (spi_data_out_r_39__N_2344[30]), 
            .\spi_data_out_r_39__N_2493[30] (spi_data_out_r_39__N_2493[30]), 
            .\spi_data_out_r_39__N_2344[29] (spi_data_out_r_39__N_2344[29]), 
            .\spi_data_out_r_39__N_2493[29] (spi_data_out_r_39__N_2493[29]), 
            .\spi_data_out_r_39__N_2344[28] (spi_data_out_r_39__N_2344[28]), 
            .\spi_data_out_r_39__N_2493[28] (spi_data_out_r_39__N_2493[28]), 
            .\spi_data_out_r_39__N_2344[27] (spi_data_out_r_39__N_2344[27]), 
            .\spi_data_out_r_39__N_2493[27] (spi_data_out_r_39__N_2493[27]), 
            .\spi_data_out_r_39__N_2344[26] (spi_data_out_r_39__N_2344[26]), 
            .\spi_data_out_r_39__N_2493[26] (spi_data_out_r_39__N_2493[26]), 
            .\spi_data_out_r_39__N_2344[25] (spi_data_out_r_39__N_2344[25]), 
            .\spi_data_out_r_39__N_2493[25] (spi_data_out_r_39__N_2493[25]), 
            .\spi_data_out_r_39__N_2344[24] (spi_data_out_r_39__N_2344[24]), 
            .\spi_data_out_r_39__N_2493[24] (spi_data_out_r_39__N_2493[24]), 
            .\spi_data_out_r_39__N_2344[23] (spi_data_out_r_39__N_2344[23]), 
            .\spi_data_out_r_39__N_2493[23] (spi_data_out_r_39__N_2493[23]), 
            .\spi_data_out_r_39__N_2344[22] (spi_data_out_r_39__N_2344[22]), 
            .\spi_data_out_r_39__N_2493[22] (spi_data_out_r_39__N_2493[22]), 
            .\spi_data_out_r_39__N_2344[21] (spi_data_out_r_39__N_2344[21]), 
            .\spi_data_out_r_39__N_2493[21] (spi_data_out_r_39__N_2493[21]), 
            .\spi_data_out_r_39__N_2344[20] (spi_data_out_r_39__N_2344[20]), 
            .\spi_data_out_r_39__N_2493[20] (spi_data_out_r_39__N_2493[20]), 
            .\spi_data_out_r_39__N_2344[19] (spi_data_out_r_39__N_2344[19]), 
            .\spi_data_out_r_39__N_2493[19] (spi_data_out_r_39__N_2493[19]), 
            .\spi_data_out_r_39__N_2344[18] (spi_data_out_r_39__N_2344[18]), 
            .\spi_data_out_r_39__N_2493[18] (spi_data_out_r_39__N_2493[18]), 
            .\spi_data_out_r_39__N_2344[17] (spi_data_out_r_39__N_2344[17]), 
            .\spi_data_out_r_39__N_2493[17] (spi_data_out_r_39__N_2493[17]), 
            .\spi_data_out_r_39__N_2344[16] (spi_data_out_r_39__N_2344[16]), 
            .\spi_data_out_r_39__N_2493[16] (spi_data_out_r_39__N_2493[16]), 
            .\spi_data_out_r_39__N_2344[15] (spi_data_out_r_39__N_2344[15]), 
            .\spi_data_out_r_39__N_2493[15] (spi_data_out_r_39__N_2493[15]), 
            .\spi_data_out_r_39__N_2344[14] (spi_data_out_r_39__N_2344[14]), 
            .\spi_data_out_r_39__N_2493[14] (spi_data_out_r_39__N_2493[14]), 
            .\spi_data_out_r_39__N_2344[13] (spi_data_out_r_39__N_2344[13]), 
            .\spi_data_out_r_39__N_2493[13] (spi_data_out_r_39__N_2493[13]), 
            .\spi_data_out_r_39__N_2344[12] (spi_data_out_r_39__N_2344[12]), 
            .\spi_data_out_r_39__N_2493[12] (spi_data_out_r_39__N_2493[12]), 
            .\spi_data_out_r_39__N_2344[11] (spi_data_out_r_39__N_2344[11]), 
            .\spi_data_out_r_39__N_2493[11] (spi_data_out_r_39__N_2493[11]), 
            .\spi_data_out_r_39__N_2344[10] (spi_data_out_r_39__N_2344[10]), 
            .\spi_data_out_r_39__N_2493[10] (spi_data_out_r_39__N_2493[10]), 
            .\spi_data_out_r_39__N_2344[9] (spi_data_out_r_39__N_2344[9]), 
            .\spi_data_out_r_39__N_2493[9] (spi_data_out_r_39__N_2493[9]), 
            .\spi_data_out_r_39__N_2344[8] (spi_data_out_r_39__N_2344[8]), 
            .\spi_data_out_r_39__N_2493[8] (spi_data_out_r_39__N_2493[8]), 
            .\spi_data_out_r_39__N_2344[7] (spi_data_out_r_39__N_2344[7]), 
            .\spi_data_out_r_39__N_2493[7] (spi_data_out_r_39__N_2493[7]), 
            .\spi_data_out_r_39__N_2344[6] (spi_data_out_r_39__N_2344[6]), 
            .\spi_data_out_r_39__N_2493[6] (spi_data_out_r_39__N_2493[6]), 
            .\spi_data_out_r_39__N_2344[5] (spi_data_out_r_39__N_2344[5]), 
            .\spi_data_out_r_39__N_2493[5] (spi_data_out_r_39__N_2493[5]), 
            .\spi_data_out_r_39__N_2344[4] (spi_data_out_r_39__N_2344[4]), 
            .\spi_data_out_r_39__N_2493[4] (spi_data_out_r_39__N_2493[4]), 
            .\spi_data_out_r_39__N_2344[3] (spi_data_out_r_39__N_2344[3]), 
            .\spi_data_out_r_39__N_2493[3] (spi_data_out_r_39__N_2493[3]), 
            .\spi_data_out_r_39__N_2344[2] (spi_data_out_r_39__N_2344[2]), 
            .\spi_data_out_r_39__N_2493[2] (spi_data_out_r_39__N_2493[2]), 
            .\spi_data_out_r_39__N_2344[1] (spi_data_out_r_39__N_2344[1]), 
            .\spi_data_out_r_39__N_2493[1] (spi_data_out_r_39__N_2493[1]), 
            .\spi_data_r[1] (spi_data_r[1]), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[3] (spi_data_r[3]), .\spi_data_r[4] (spi_data_r[4]), 
            .\spi_data_r[5] (spi_data_r[5]), .\spi_data_r[6] (spi_data_r[6]), 
            .\spi_data_r[7] (spi_data_r[7]), .\spi_data_r[8] (spi_data_r[8]), 
            .\spi_data_r[9] (spi_data_r[9]), .\spi_data_r[10] (spi_data_r[10]), 
            .\spi_data_r[11] (spi_data_r[11]), .\spi_data_r[12] (spi_data_r[12]), 
            .\spi_data_r[13] (spi_data_r[13]), .\spi_data_r[14] (spi_data_r[14]), 
            .\spi_data_r[15] (spi_data_r[15]), .\spi_data_r[16] (spi_data_r[16]), 
            .\spi_data_r[17] (spi_data_r[17]), .\spi_data_r[18] (spi_data_r[18]), 
            .\spi_data_r[19] (spi_data_r[19]), .\spi_data_r[20] (spi_data_r[20]), 
            .\spi_data_r[21] (spi_data_r[21]), .\spi_data_r[22] (spi_data_r[22]), 
            .\spi_data_r[23] (spi_data_r[23]), .\spi_data_r[24] (spi_data_r[24]), 
            .\spi_data_r[25] (spi_data_r[25]), .\spi_data_r[26] (spi_data_r[26]), 
            .\spi_data_r[27] (spi_data_r[27]), .\spi_data_r[28] (spi_data_r[28]), 
            .\spi_data_r[29] (spi_data_r[29]), .\spi_data_r[30] (spi_data_r[30]), 
            .\spi_data_r[31] (spi_data_r[31]), .resetn_c(resetn_c), .n1(n1_adj_7667)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(263[3] 283[2])
    \peizo_elliptec(DEV_ID=7,UART_ADDRESS_WIDTH=4)  u_peizo_elliptec (.mode(mode_adj_7729), 
            .clk(clk), .clk_enable_32(clk_enable_32), .n30185(n30185), 
            .\spi_data_r[0] (spi_data_r[0]), .n28(n28), .n29594(n29594), 
            .uart_slot_en({uart_slot_en}), .n30118(n30118), .n6(n6), .n29944(n29944), 
            .n29943(n29943), .\spi_cmd_r[0] (spi_cmd_r[0]), .spi_addr_r({spi_addr_r}), 
            .n30138(n30138), .\spi_cmd_r[2] (spi_cmd_r[2]), .n30023(n30023), 
            .n26107(n26107), .n30090(n30090), .n29481(n29481), .n25941(n25941), 
            .n25923(n25923), .n30062(n30062), .n30087(n30087), .pin_io_out_55(pin_io_out_55), 
            .n28358(n28358), .pin_io_out_40(pin_io_out_40), .n30122(n30122), 
            .n24700(n24700), .n23248(n23248), .n10696(n10696), .tx_N_6586(tx_N_6586), 
            .n25358(n25358), .n30083(n30083), .mode_adj_656(mode_adj_7727), 
            .C_8_c(C_8_c), .n30064(n30064), .n30155(n30155), .n26091(n26091), 
            .n30214(n30214), .n28402(n28402), .n30094(n30094), .n28486(n28486), 
            .n18440(n18440), .n26113(n26113), .n26119(n26119), .n30095(n30095), 
            .pin_io_out_25(pin_io_out_25), .mode_adj_657(mode_adj_7725), 
            .n30043(n30043), .n4(n4_adj_7733), .pin_io_out_6(pin_io_out_6), 
            .mode_adj_658(mode), .mode_adj_659(mode_adj_7724), .pin_io_out_5(pin_io_out_5), 
            .n30120(n30120), .n23409(n23409), .n26089(n26089), .n25739(n25739), 
            .n25741(n25741)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(591[3] 611[2])
    \intrpt_ctrl(DEV_ID=4)  \intrpt_ins_4..u_intrpt_ctrl  (.clk(clk), .n30185(n30185), 
            .\pin_intrpt[12] (pin_intrpt[12]), .intrpt_out_c_4(intrpt_out_c_4), 
            .intrpt_out_N_2926(intrpt_out_N_2926), .n31069(n31069), .\spi_data_out_r_39__N_2863[0] (spi_data_out_r_39__N_2863[0]), 
            .clear_intrpt(clear_intrpt_adj_7664), .clear_intrpt_N_2930(clear_intrpt_N_2930), 
            .\spi_data_out_r_39__N_2863[2] (spi_data_out_r_39__N_2863[2]), 
            .\pin_intrpt[14] (pin_intrpt[14]), .\spi_data_out_r_39__N_2863[1] (spi_data_out_r_39__N_2863[1]), 
            .\pin_intrpt[13] (pin_intrpt[13])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(294[3] 315[2])
    \intrpt_ctrl(DEV_ID=6)  \intrpt_ins_6..u_intrpt_ctrl  (.clk(clk), .n30185(n30185), 
            .\spi_data_out_r_39__N_3005[0] (spi_data_out_r_39__N_3005[0]), 
            .\pin_intrpt[18] (pin_intrpt[18]), .intrpt_out_c_6(intrpt_out_c_6), 
            .intrpt_out_N_3068(intrpt_out_N_3068), .n31069(n31069), .\spi_data_out_r_39__N_3005[2] (spi_data_out_r_39__N_3005[2]), 
            .\pin_intrpt[20] (pin_intrpt[20]), .\spi_data_out_r_39__N_3005[1] (spi_data_out_r_39__N_3005[1]), 
            .\pin_intrpt[19] (pin_intrpt[19]), .clear_intrpt(clear_intrpt_adj_7666), 
            .clear_intrpt_N_3072(clear_intrpt_N_3072)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(294[3] 315[2])
    \status_led(DEV_ID=9)  u_status_led (.clk(clk), .clk_enable_595(clk_enable_595), 
            .n30185(n30185), .\spi_data_r[0] (spi_data_r[0]), .\spi_data_out_r_39__N_770[0] (spi_data_out_r_39__N_770[0]), 
            .GND_net(GND_net), .n30039(n30039), .n12435(n12435), .spi_data_out_r_39__N_810(spi_data_out_r_39__N_810), 
            .n12467(n12467), .\status_cntr[11] (status_cntr[11]), .\status_cntr[12] (status_cntr[12]), 
            .n18654(n18654), .EM_STOP(EM_STOP), .led_sw_c(led_sw_c), .clk_enable_227(clk_enable_227), 
            .n25212(n25212), .n4(n4), .\spi_data_r[11] (spi_data_r[11]), 
            .\spi_data_r[10] (spi_data_r[10]), .\spi_data_r[9] (spi_data_r[9]), 
            .\spi_data_r[8] (spi_data_r[8]), .\spi_data_r[7] (spi_data_r[7]), 
            .\spi_data_r[6] (spi_data_r[6]), .\spi_data_r[5] (spi_data_r[5]), 
            .\spi_data_r[4] (spi_data_r[4]), .\spi_data_r[3] (spi_data_r[3]), 
            .\spi_data_r[2] (spi_data_r[2]), .\spi_data_r[1] (spi_data_r[1]), 
            .pwm(pwm), .resetn_c(resetn_c), .n28562(n28562), .n57(n57), 
            .n6651(n6651), .pwm_duty_3({pwm_duty_3_adj_8331}), .n21(n21_adj_7737), 
            .n19(n19_adj_7736), .n20(n20), .n6649(n6649), .pwm_N_898(pwm_N_898), 
            .n22554(n22554), .pwm_N_896(pwm_N_896), .n6747(n6747), .pwm_duty_1({pwm_duty_1_adj_8329}), 
            .n30020(n30020), .n20647(n20647), .n6590(n6590), .pwm_duty_2({pwm_duty_2_adj_8330}), 
            .n30102(n30102), .n29997(n29997), .\spi_cmd[2] (spi_cmd[2]), 
            .n27095(n27095)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(219[3] 236[2])
    LUT4 i23843_4_lut_else_4_lut (.A(cs_c_4), .B(cs_c_3), .C(cs_c_2), 
         .D(cs_c_0), .Z(n30218)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i23843_4_lut_else_4_lut.init = 16'h0001;
    pll __ (.clk_in_c(clk_in_c), .clk_100k(clk_100k), .clk_1MHz(clk_1MHz), 
        .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(140[5:100])
    TSALL TSALL_INST (.TSALL(GND_net));
    LUT4 m1_lut (.Z(n31069)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    GSR GSR_INST (.GSR(resetn_c));
    pwm_controller \pwm_ins_0..pwm_controller_ins  (.\pwm_out[0] (pwm_out[0]), 
            .clk(clk), .clk_enable_15(clk_enable_15), .n2109(n2109), .clk_enable_263(clk_enable_263), 
            .n30185(n30185), .\spi_data_r[0] (spi_data_r[0]), .clk_enable_638(clk_enable_638), 
            .\spi_data_r[11] (spi_data_r[11]), .\spi_data_r[10] (spi_data_r[10]), 
            .\spi_data_r[9] (spi_data_r[9]), .\spi_data_r[8] (spi_data_r[8]), 
            .\spi_data_r[7] (spi_data_r[7]), .\spi_data_r[6] (spi_data_r[6]), 
            .\spi_data_r[5] (spi_data_r[5]), .\spi_data_r[4] (spi_data_r[4]), 
            .\spi_data_r[3] (spi_data_r[3]), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[1] (spi_data_r[1]), .GND_net(GND_net), .pwm_out_N_3153(pwm_out_N_3153), 
            .pwm_out_N_3169(pwm_out_N_3169), .resetn_c(resetn_c)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(327[5] 339[4])
    \quad_decoder(DEV_ID=4)  \quad_ins_4..u_quad_decoder  (.quad_count({quad_count_adj_7892}), 
            .clk(clk), .n30185(n30185), .\quad_a[4] (quad_a[4]), .\quad_b[4] (quad_b[4]), 
            .\spi_data_out_r_39__N_1874[0] (spi_data_out_r_39__N_1874[0]), 
            .\spi_data_out_r_39__N_2023[0] (spi_data_out_r_39__N_2023[0]), 
            .quad_buffer({quad_buffer_adj_7893}), .\pin_intrpt[14] (pin_intrpt[14]), 
            .clk_enable_683(clk_enable_683), .\spi_data_r[0] (spi_data_r[0]), 
            .quad_homing({quad_homing_adj_7891}), .clk_enable_684(clk_enable_684), 
            .spi_data_out_r_39__N_1914(spi_data_out_r_39__N_1914), .spi_data_out_r_39__N_2103(spi_data_out_r_39__N_2103), 
            .quad_set_valid_N_2098(quad_set_valid_N_2098), .\spi_data_out_r_39__N_1874[31] (spi_data_out_r_39__N_1874[31]), 
            .\spi_data_out_r_39__N_2023[31] (spi_data_out_r_39__N_2023[31]), 
            .\spi_data_out_r_39__N_1874[30] (spi_data_out_r_39__N_1874[30]), 
            .\spi_data_out_r_39__N_2023[30] (spi_data_out_r_39__N_2023[30]), 
            .\spi_data_out_r_39__N_1874[29] (spi_data_out_r_39__N_1874[29]), 
            .\spi_data_out_r_39__N_2023[29] (spi_data_out_r_39__N_2023[29]), 
            .\spi_data_out_r_39__N_1874[28] (spi_data_out_r_39__N_1874[28]), 
            .\spi_data_out_r_39__N_2023[28] (spi_data_out_r_39__N_2023[28]), 
            .\spi_data_out_r_39__N_1874[27] (spi_data_out_r_39__N_1874[27]), 
            .\spi_data_out_r_39__N_2023[27] (spi_data_out_r_39__N_2023[27]), 
            .\spi_data_out_r_39__N_1874[26] (spi_data_out_r_39__N_1874[26]), 
            .\spi_data_out_r_39__N_2023[26] (spi_data_out_r_39__N_2023[26]), 
            .\spi_data_out_r_39__N_1874[25] (spi_data_out_r_39__N_1874[25]), 
            .\spi_data_out_r_39__N_2023[25] (spi_data_out_r_39__N_2023[25]), 
            .\spi_data_out_r_39__N_1874[24] (spi_data_out_r_39__N_1874[24]), 
            .\spi_data_out_r_39__N_2023[24] (spi_data_out_r_39__N_2023[24]), 
            .\spi_data_out_r_39__N_1874[23] (spi_data_out_r_39__N_1874[23]), 
            .\spi_data_out_r_39__N_2023[23] (spi_data_out_r_39__N_2023[23]), 
            .\spi_data_out_r_39__N_1874[22] (spi_data_out_r_39__N_1874[22]), 
            .\spi_data_out_r_39__N_2023[22] (spi_data_out_r_39__N_2023[22]), 
            .\spi_data_out_r_39__N_1874[21] (spi_data_out_r_39__N_1874[21]), 
            .\spi_data_out_r_39__N_2023[21] (spi_data_out_r_39__N_2023[21]), 
            .\spi_data_out_r_39__N_1874[20] (spi_data_out_r_39__N_1874[20]), 
            .\spi_data_out_r_39__N_2023[20] (spi_data_out_r_39__N_2023[20]), 
            .\spi_data_out_r_39__N_1874[19] (spi_data_out_r_39__N_1874[19]), 
            .\spi_data_out_r_39__N_2023[19] (spi_data_out_r_39__N_2023[19]), 
            .\spi_data_out_r_39__N_1874[18] (spi_data_out_r_39__N_1874[18]), 
            .\spi_data_out_r_39__N_2023[18] (spi_data_out_r_39__N_2023[18]), 
            .\spi_data_out_r_39__N_1874[17] (spi_data_out_r_39__N_1874[17]), 
            .\spi_data_out_r_39__N_2023[17] (spi_data_out_r_39__N_2023[17]), 
            .\spi_data_out_r_39__N_1874[16] (spi_data_out_r_39__N_1874[16]), 
            .\spi_data_out_r_39__N_2023[16] (spi_data_out_r_39__N_2023[16]), 
            .\spi_data_out_r_39__N_1874[15] (spi_data_out_r_39__N_1874[15]), 
            .\spi_data_out_r_39__N_2023[15] (spi_data_out_r_39__N_2023[15]), 
            .\spi_data_out_r_39__N_1874[14] (spi_data_out_r_39__N_1874[14]), 
            .\spi_data_out_r_39__N_2023[14] (spi_data_out_r_39__N_2023[14]), 
            .\spi_data_out_r_39__N_1874[13] (spi_data_out_r_39__N_1874[13]), 
            .\spi_data_out_r_39__N_2023[13] (spi_data_out_r_39__N_2023[13]), 
            .\spi_data_out_r_39__N_1874[12] (spi_data_out_r_39__N_1874[12]), 
            .\spi_data_out_r_39__N_2023[12] (spi_data_out_r_39__N_2023[12]), 
            .\spi_data_out_r_39__N_1874[11] (spi_data_out_r_39__N_1874[11]), 
            .\spi_data_out_r_39__N_2023[11] (spi_data_out_r_39__N_2023[11]), 
            .\spi_data_out_r_39__N_1874[10] (spi_data_out_r_39__N_1874[10]), 
            .\spi_data_out_r_39__N_2023[10] (spi_data_out_r_39__N_2023[10]), 
            .\spi_data_out_r_39__N_1874[9] (spi_data_out_r_39__N_1874[9]), 
            .\spi_data_out_r_39__N_2023[9] (spi_data_out_r_39__N_2023[9]), 
            .\spi_data_out_r_39__N_1874[8] (spi_data_out_r_39__N_1874[8]), 
            .\spi_data_out_r_39__N_2023[8] (spi_data_out_r_39__N_2023[8]), 
            .\spi_data_out_r_39__N_1874[7] (spi_data_out_r_39__N_1874[7]), 
            .\spi_data_out_r_39__N_2023[7] (spi_data_out_r_39__N_2023[7]), 
            .\spi_data_out_r_39__N_1874[6] (spi_data_out_r_39__N_1874[6]), 
            .\spi_data_out_r_39__N_2023[6] (spi_data_out_r_39__N_2023[6]), 
            .\spi_data_out_r_39__N_1874[5] (spi_data_out_r_39__N_1874[5]), 
            .\spi_data_out_r_39__N_2023[5] (spi_data_out_r_39__N_2023[5]), 
            .\spi_data_out_r_39__N_1874[4] (spi_data_out_r_39__N_1874[4]), 
            .\spi_data_out_r_39__N_2023[4] (spi_data_out_r_39__N_2023[4]), 
            .\spi_data_out_r_39__N_1874[3] (spi_data_out_r_39__N_1874[3]), 
            .\spi_data_out_r_39__N_2023[3] (spi_data_out_r_39__N_2023[3]), 
            .\spi_data_out_r_39__N_1874[2] (spi_data_out_r_39__N_1874[2]), 
            .\spi_data_out_r_39__N_2023[2] (spi_data_out_r_39__N_2023[2]), 
            .\spi_data_out_r_39__N_1874[1] (spi_data_out_r_39__N_1874[1]), 
            .\spi_data_out_r_39__N_2023[1] (spi_data_out_r_39__N_2023[1]), 
            .n1(n1_adj_7712), .\spi_data_r[1] (spi_data_r[1]), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[3] (spi_data_r[3]), .\spi_data_r[4] (spi_data_r[4]), 
            .\spi_data_r[5] (spi_data_r[5]), .\spi_data_r[6] (spi_data_r[6]), 
            .\spi_data_r[7] (spi_data_r[7]), .\spi_data_r[8] (spi_data_r[8]), 
            .\spi_data_r[9] (spi_data_r[9]), .\spi_data_r[10] (spi_data_r[10]), 
            .\spi_data_r[11] (spi_data_r[11]), .\spi_data_r[12] (spi_data_r[12]), 
            .\spi_data_r[13] (spi_data_r[13]), .\spi_data_r[14] (spi_data_r[14]), 
            .\spi_data_r[15] (spi_data_r[15]), .\spi_data_r[16] (spi_data_r[16]), 
            .\spi_data_r[17] (spi_data_r[17]), .\spi_data_r[18] (spi_data_r[18]), 
            .\spi_data_r[19] (spi_data_r[19]), .\spi_data_r[20] (spi_data_r[20]), 
            .\spi_data_r[21] (spi_data_r[21]), .\spi_data_r[22] (spi_data_r[22]), 
            .\spi_data_r[23] (spi_data_r[23]), .\spi_data_r[24] (spi_data_r[24]), 
            .\spi_data_r[25] (spi_data_r[25]), .\spi_data_r[26] (spi_data_r[26]), 
            .\spi_data_r[27] (spi_data_r[27]), .\spi_data_r[28] (spi_data_r[28]), 
            .\spi_data_r[29] (spi_data_r[29]), .\spi_data_r[30] (spi_data_r[30]), 
            .\spi_data_r[31] (spi_data_r[31]), .GND_net(GND_net), .resetn_c(resetn_c)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(263[3] 283[2])
    PFUMX i24393 (.BLUT(n30218), .ALUT(n30219), .C0(FLASH_CS_c), .Z(n30220));
    \rs232(DEV_ID=4,UART_ADDRESS_WIDTH=4)  u_rs232 (.n28340(n28340), .n24066(n24066), 
            .n28328(n28328), .quad_set_valid_N_2333(quad_set_valid_N_2333), 
            .spi_addr_r({spi_addr_r}), .n30214(n30214), .n25643(n25643), 
            .n30210(n30210), .mode(mode_adj_7727), .clk(clk), .clk_enable_253(clk_enable_253), 
            .n30185(n30185), .\spi_data_r[0] (spi_data_r[0]), .\spi_cmd_r[0] (spi_cmd_r[0]), 
            .n26107(n26107), .n26621(n26621), .n26207(n26207), .n30071(n30071), 
            .\spi_cmd_r[5] (spi_cmd_r[5]), .n28476(n28476), .n26819(n26819), 
            .n30144(n30144), .n26821(n26821), .\spi_cmd_r[3] (spi_cmd_r[3]), 
            .n30155(n30155), .n28260(n28260), .n30044(n30044), .n25941(n25941), 
            .n18440(n18440), .n30213(n30213), .n25979(n25979), .resetn_c(resetn_c), 
            .n30122(n30122), .\uart_slot_en[0] (uart_slot_en[0]), .\uart_slot_en[2] (uart_slot_en[2]), 
            .\uart_slot_en[1] (uart_slot_en[1]), .TX_IN_N_6565(TX_IN_N_6565), 
            .n25739(n25739), .UC_TXD0_c(UC_TXD0_c), .n30180(n30180), .n7164(n7164), 
            .n26633(n26633), .n23916(n23916), .n23526(n23526), .n30004(n30004), 
            .n26947(n26947), .\spi_cmd_r[2] (spi_cmd_r[2]), .n30199(n30199), 
            .n30031(n30031)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(541[3] 561[2])
    \stepper(DEV_ID=2,UART_ADDRESS_WIDTH=4)  \stepper_ins_2..u_stepper  (.clk(clk), 
            .clk_1MHz(clk_1MHz), .n30185(n30185), .GND_net(GND_net), .pin_io_c_28(pin_io_c_28), 
            .reset_r(reset_r_adj_7676), .clk_enable_23(clk_enable_23), .n29996(n29996), 
            .resetn_c(resetn_c), .n30110(n30110), .spi_data_out_r_39__N_4511({spi_data_out_r_39__N_4511}), 
            .clk_enable_686(clk_enable_686), .\spi_data_r[0] (spi_data_r[0]), 
            .n47(n47_adj_7731), .spi_data_out_r_39__N_4551(spi_data_out_r_39__N_4551), 
            .spi_data_out_r_39__N_4848(spi_data_out_r_39__N_4848), .digital_output_r(digital_output_r_adj_7677), 
            .clk_enable_259(clk_enable_259), .n28556(n28556), .\quad_homing[0] (quad_homing_adj_7815[0]), 
            .pin_io_c_24(pin_io_c_24), .n25881(n25881), .\spi_data_r[1] (spi_data_r[1]), 
            .\mode[2] (n31091[2]), .\spi_data_r[2] (spi_data_r[2]), .NSL(NSL_adj_7678), 
            .n5(n5_adj_7726), .UC_TXD0_c(UC_TXD0_c), .OW_ID_N_4804(OW_ID_N_4804), 
            .n9(n9_adj_7674), .\uart_slot_en[0] (uart_slot_en[0]), .\uart_slot_en[1] (uart_slot_en[1]), 
            .pin_io_out_29(pin_io_out_29), .\quad_b[2] (quad_b[2]), .\quad_a[2] (quad_a[2]), 
            .pin_io_c_23(pin_io_c_23), .\pin_intrpt[7] (pin_intrpt[7]), 
            .n30095(n30095), .OW_ID_N_4810(OW_ID_N_4810), .pin_io_c_22(pin_io_c_22), 
            .\pin_intrpt[6] (pin_intrpt[6]), .\pin_intrpt[8] (pin_intrpt[8]), 
            .n7273(n7273), .ENC_O_N_4812(ENC_O_N_4812)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(354[3] 397[2])
    \quad_decoder(DEV_ID=5)  \quad_ins_5..u_quad_decoder  (.quad_homing({quad_homing_adj_7929}), 
            .clk(clk), .clk_enable_388(clk_enable_388), .n30185(n30185), 
            .\spi_data_r[0] (spi_data_r[0]), .quad_count({quad_count_adj_7930}), 
            .\quad_b[5] (quad_b[5]), .\spi_data_out_r_39__N_2109[0] (spi_data_out_r_39__N_2109[0]), 
            .\spi_data_out_r_39__N_2258[0] (spi_data_out_r_39__N_2258[0]), 
            .quad_buffer({quad_buffer_adj_7931}), .\pin_intrpt[17] (pin_intrpt[17]), 
            .GND_net(GND_net), .clk_enable_315(clk_enable_315), .\quad_a[5] (quad_a[5]), 
            .spi_data_out_r_39__N_2149(spi_data_out_r_39__N_2149), .spi_data_out_r_39__N_2338(spi_data_out_r_39__N_2338), 
            .quad_set_valid_N_2333(quad_set_valid_N_2333), .\spi_data_r[31] (spi_data_r[31]), 
            .\spi_data_r[30] (spi_data_r[30]), .\spi_data_r[29] (spi_data_r[29]), 
            .\spi_data_r[28] (spi_data_r[28]), .\spi_data_r[27] (spi_data_r[27]), 
            .\spi_data_r[26] (spi_data_r[26]), .\spi_data_r[25] (spi_data_r[25]), 
            .\spi_data_r[24] (spi_data_r[24]), .\spi_data_r[23] (spi_data_r[23]), 
            .\spi_data_r[22] (spi_data_r[22]), .\spi_data_r[21] (spi_data_r[21]), 
            .\spi_data_r[20] (spi_data_r[20]), .\spi_data_r[19] (spi_data_r[19]), 
            .\spi_data_r[18] (spi_data_r[18]), .\spi_data_r[17] (spi_data_r[17]), 
            .\spi_data_r[16] (spi_data_r[16]), .\spi_data_r[15] (spi_data_r[15]), 
            .\spi_data_r[14] (spi_data_r[14]), .\spi_data_r[13] (spi_data_r[13]), 
            .\spi_data_r[12] (spi_data_r[12]), .\spi_data_r[11] (spi_data_r[11]), 
            .\spi_data_r[10] (spi_data_r[10]), .\spi_data_r[9] (spi_data_r[9]), 
            .\spi_data_r[8] (spi_data_r[8]), .\spi_data_r[7] (spi_data_r[7]), 
            .\spi_data_r[6] (spi_data_r[6]), .\spi_data_r[5] (spi_data_r[5]), 
            .\spi_data_r[4] (spi_data_r[4]), .\spi_data_r[3] (spi_data_r[3]), 
            .\spi_data_r[2] (spi_data_r[2]), .\spi_data_r[1] (spi_data_r[1]), 
            .\spi_data_out_r_39__N_2109[31] (spi_data_out_r_39__N_2109[31]), 
            .\spi_data_out_r_39__N_2258[31] (spi_data_out_r_39__N_2258[31]), 
            .\spi_data_out_r_39__N_2109[30] (spi_data_out_r_39__N_2109[30]), 
            .\spi_data_out_r_39__N_2258[30] (spi_data_out_r_39__N_2258[30]), 
            .\spi_data_out_r_39__N_2109[29] (spi_data_out_r_39__N_2109[29]), 
            .\spi_data_out_r_39__N_2258[29] (spi_data_out_r_39__N_2258[29]), 
            .\spi_data_out_r_39__N_2109[28] (spi_data_out_r_39__N_2109[28]), 
            .\spi_data_out_r_39__N_2258[28] (spi_data_out_r_39__N_2258[28]), 
            .\spi_data_out_r_39__N_2109[27] (spi_data_out_r_39__N_2109[27]), 
            .\spi_data_out_r_39__N_2258[27] (spi_data_out_r_39__N_2258[27]), 
            .\spi_data_out_r_39__N_2109[26] (spi_data_out_r_39__N_2109[26]), 
            .\spi_data_out_r_39__N_2258[26] (spi_data_out_r_39__N_2258[26]), 
            .\spi_data_out_r_39__N_2109[25] (spi_data_out_r_39__N_2109[25]), 
            .\spi_data_out_r_39__N_2258[25] (spi_data_out_r_39__N_2258[25]), 
            .\spi_data_out_r_39__N_2109[24] (spi_data_out_r_39__N_2109[24]), 
            .\spi_data_out_r_39__N_2258[24] (spi_data_out_r_39__N_2258[24]), 
            .\spi_data_out_r_39__N_2109[23] (spi_data_out_r_39__N_2109[23]), 
            .\spi_data_out_r_39__N_2258[23] (spi_data_out_r_39__N_2258[23]), 
            .\spi_data_out_r_39__N_2109[22] (spi_data_out_r_39__N_2109[22]), 
            .\spi_data_out_r_39__N_2258[22] (spi_data_out_r_39__N_2258[22]), 
            .\spi_data_out_r_39__N_2109[21] (spi_data_out_r_39__N_2109[21]), 
            .\spi_data_out_r_39__N_2258[21] (spi_data_out_r_39__N_2258[21]), 
            .\spi_data_out_r_39__N_2109[20] (spi_data_out_r_39__N_2109[20]), 
            .\spi_data_out_r_39__N_2258[20] (spi_data_out_r_39__N_2258[20]), 
            .\spi_data_out_r_39__N_2109[19] (spi_data_out_r_39__N_2109[19]), 
            .\spi_data_out_r_39__N_2258[19] (spi_data_out_r_39__N_2258[19]), 
            .\spi_data_out_r_39__N_2109[18] (spi_data_out_r_39__N_2109[18]), 
            .\spi_data_out_r_39__N_2258[18] (spi_data_out_r_39__N_2258[18]), 
            .\spi_data_out_r_39__N_2109[17] (spi_data_out_r_39__N_2109[17]), 
            .\spi_data_out_r_39__N_2258[17] (spi_data_out_r_39__N_2258[17]), 
            .\spi_data_out_r_39__N_2109[16] (spi_data_out_r_39__N_2109[16]), 
            .\spi_data_out_r_39__N_2258[16] (spi_data_out_r_39__N_2258[16]), 
            .\spi_data_out_r_39__N_2109[15] (spi_data_out_r_39__N_2109[15]), 
            .\spi_data_out_r_39__N_2258[15] (spi_data_out_r_39__N_2258[15]), 
            .\spi_data_out_r_39__N_2109[14] (spi_data_out_r_39__N_2109[14]), 
            .\spi_data_out_r_39__N_2258[14] (spi_data_out_r_39__N_2258[14]), 
            .\spi_data_out_r_39__N_2109[13] (spi_data_out_r_39__N_2109[13]), 
            .\spi_data_out_r_39__N_2258[13] (spi_data_out_r_39__N_2258[13]), 
            .\spi_data_out_r_39__N_2109[12] (spi_data_out_r_39__N_2109[12]), 
            .\spi_data_out_r_39__N_2258[12] (spi_data_out_r_39__N_2258[12]), 
            .\spi_data_out_r_39__N_2109[11] (spi_data_out_r_39__N_2109[11]), 
            .\spi_data_out_r_39__N_2258[11] (spi_data_out_r_39__N_2258[11]), 
            .\spi_data_out_r_39__N_2109[10] (spi_data_out_r_39__N_2109[10]), 
            .\spi_data_out_r_39__N_2258[10] (spi_data_out_r_39__N_2258[10]), 
            .\spi_data_out_r_39__N_2109[9] (spi_data_out_r_39__N_2109[9]), 
            .\spi_data_out_r_39__N_2258[9] (spi_data_out_r_39__N_2258[9]), 
            .\spi_data_out_r_39__N_2109[8] (spi_data_out_r_39__N_2109[8]), 
            .\spi_data_out_r_39__N_2258[8] (spi_data_out_r_39__N_2258[8]), 
            .\spi_data_out_r_39__N_2109[7] (spi_data_out_r_39__N_2109[7]), 
            .\spi_data_out_r_39__N_2258[7] (spi_data_out_r_39__N_2258[7]), 
            .\spi_data_out_r_39__N_2109[6] (spi_data_out_r_39__N_2109[6]), 
            .\spi_data_out_r_39__N_2258[6] (spi_data_out_r_39__N_2258[6]), 
            .\spi_data_out_r_39__N_2109[5] (spi_data_out_r_39__N_2109[5]), 
            .\spi_data_out_r_39__N_2258[5] (spi_data_out_r_39__N_2258[5]), 
            .\spi_data_out_r_39__N_2109[4] (spi_data_out_r_39__N_2109[4]), 
            .\spi_data_out_r_39__N_2258[4] (spi_data_out_r_39__N_2258[4]), 
            .\spi_data_out_r_39__N_2109[3] (spi_data_out_r_39__N_2109[3]), 
            .\spi_data_out_r_39__N_2258[3] (spi_data_out_r_39__N_2258[3]), 
            .\spi_data_out_r_39__N_2109[2] (spi_data_out_r_39__N_2109[2]), 
            .\spi_data_out_r_39__N_2258[2] (spi_data_out_r_39__N_2258[2]), 
            .\spi_data_out_r_39__N_2109[1] (spi_data_out_r_39__N_2109[1]), 
            .\spi_data_out_r_39__N_2258[1] (spi_data_out_r_39__N_2258[1]), 
            .resetn_c(resetn_c), .n1(n1_adj_7669)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(263[3] 283[2])
    \servo(UART_ADDRESS_WIDTH=4)  \servo_ins_0..u_servo  (.pin_io_out_2(pin_io_out_2), 
            .pin_io_out_1(pin_io_out_1), .n30043(n30043), .mode(mode), 
            .\pin_intrpt[0] (pin_intrpt[0]), .clk(clk), .clk_enable_232(clk_enable_232), 
            .n30185(n30185), .\spi_data_r[0] (spi_data_r[0]), .Phase_r(Phase_r), 
            .clk_enable_234(clk_enable_234), .pin_io_out_9(pin_io_out_9), 
            .\quad_b[0] (quad_b[0]), .mode_adj_655({n31089}), .\spi_cmd_r[2] (spi_cmd_r[2]), 
            .\spi_cmd_r[0] (spi_cmd_r[0]), .n23732(n23732), .pin_io_out_8(pin_io_out_8), 
            .\quad_a[0] (quad_a[0]), .\uart_slot_en[3] (uart_slot_en[3]), 
            .\uart_slot_en[0] (uart_slot_en[0]), .n8(n8), .pin_io_out_3(pin_io_out_3), 
            .\pin_intrpt[1] (pin_intrpt[1])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(408[3] 443[2])
    \otm_dac(DEV_ID=3)  u_otm_dac (.clk(clk), .clk_enable_255(clk_enable_255), 
            .n30185(n30185), .\spi_data_r[0] (spi_data_r[0]), .mode(mode_adj_7728), 
            .clk_enable_260(clk_enable_260), .NSL(NSL_adj_7681), .n30082(n30082), 
            .n7167(n7167)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(566[3] 584[2])
    \stepper(DEV_ID=5,UART_ADDRESS_WIDTH=4)  \stepper_ins_5..u_stepper  (.clk_1MHz(clk_1MHz), 
            .n30185(n30185), .clk(clk), .reset_r(reset_r_adj_7717), .clk_enable_38(clk_enable_38), 
            .n29994(n29994), .clk_enable_627(clk_enable_627), .\spi_data_r[0] (spi_data_r[0]), 
            .GND_net(GND_net), .pin_io_c_58(pin_io_c_58), .n30149(n30149), 
            .spi_data_out_r_39__N_5540({spi_data_out_r_39__N_5540}), .resetn_c(resetn_c), 
            .digital_output_r(digital_output_r_adj_7718), .clk_enable_242(clk_enable_242), 
            .n28551(n28551), .spi_data_out_r_39__N_5580(spi_data_out_r_39__N_5580), 
            .spi_data_out_r_39__N_5877(spi_data_out_r_39__N_5877), .\spi_data_r[1] (spi_data_r[1]), 
            .\spi_data_r[2] (spi_data_r[2]), .n47(n47_adj_7716), .NSL(NSL_adj_7719), 
            .\uart_slot_en[2] (uart_slot_en[2]), .\uart_slot_en[3] (uart_slot_en[3]), 
            .n10696(n10696), .\quad_homing[0] (quad_homing_adj_7929[0]), 
            .pin_io_c_54(pin_io_c_54), .n25885(n25885), .pin_io_out_59(pin_io_out_59), 
            .\quad_b[5] (quad_b[5]), .UC_TXD0_c(UC_TXD0_c), .OW_ID_N_5833(OW_ID_N_5833), 
            .OW_ID_N_5839(OW_ID_N_5839), .n30049(n30049), .\uart_slot_en[0] (uart_slot_en[0]), 
            .\quad_a[5] (quad_a[5]), .n30047(n30047), .n30087(n30087), 
            .\pin_intrpt[17] (pin_intrpt[17]), .n7262(n7262), .pin_io_c_52(pin_io_c_52), 
            .\pin_intrpt[15] (pin_intrpt[15]), .pin_io_c_53(pin_io_c_53), 
            .\pin_intrpt[16] (pin_intrpt[16]), .ENC_O_N_5841(ENC_O_N_5841)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(354[3] 397[2])
    \io(UART_ADDRESS_WIDTH=4)  \io_ins_0..u_io  (.pwm_out_1(pwm_out_1), .clk_100k(clk_100k), 
            .clk_100k_enable_1(clk_100k_enable_1), .n2193(n2193), .clk(clk), 
            .clk_enable_695(clk_enable_695), .n30185(n30185), .\spi_data_r[0] (spi_data_r[0]), 
            .mode(mode_adj_7724), .clk_enable_235(clk_enable_235), .\spi_data_r[1] (spi_data_r[1]), 
            .\spi_data_r[3] (spi_data_r[3]), .\spi_data_r[4] (spi_data_r[4]), 
            .\spi_data_r[7] (spi_data_r[7]), .\spi_data_r[8] (spi_data_r[8]), 
            .\spi_data_r[9] (spi_data_r[9]), .\spi_data_r[10] (spi_data_r[10]), 
            .\spi_data_r[11] (spi_data_r[11]), .GND_net(GND_net), .pwm_out_1_N_6306(pwm_out_1_N_6306), 
            .clk_enable_959(clk_enable_959), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[5] (spi_data_r[5]), .\spi_data_r[6] (spi_data_r[6]), 
            .n18(n18), .resetn_c(resetn_c)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(454[3] 486[2])
    \stepper(UART_ADDRESS_WIDTH=4)  \stepper_ins_0..u_stepper  (.GND_net(GND_net), 
            .clk(clk), .\spi_addr_r[0] (spi_addr_r[0]), .n30070(n30070), 
            .n23526(n23526), .n30035(n30035), .n29990(n29990), .clk_1MHz(clk_1MHz), 
            .n30185(n30185), .resetn_c(resetn_c), .n30129(n30129), .spi_data_out_r_39__N_3825({spi_data_out_r_39__N_3825}), 
            .pin_io_out_8(pin_io_out_8), .spi_data_out_r_39__N_3865(spi_data_out_r_39__N_3865), 
            .mode_adj_654({n31089}), .clk_enable_761(clk_enable_761), .\spi_data_r[0] (spi_data_r[0]), 
            .n30175(n30175), .n30058(n30058), .digital_output_r(digital_output_r), 
            .n28547(n28547), .n47(n47_adj_7732), .\spi_addr_r[1] (spi_addr_r[1]), 
            .n26957(n26957), .n23537(n23537), .n20647(n20647), .n23978(n23978), 
            .\spi_cmd_r[2] (spi_cmd_r[2]), .\spi_cmd_r[8] (spi_cmd_r[8]), 
            .\spi_cmd_r[10] (spi_cmd_r[10]), .\spi_cmd_r[6] (spi_cmd_r[6]), 
            .\spi_cmd_r[7] (spi_cmd_r[7]), .\spi_cmd_r[12] (spi_cmd_r[12]), 
            .\spi_cmd_r[15] (spi_cmd_r[15]), .n30134(n30134), .n30125(n30125), 
            .mode(mode), .n23609(n23609), .n30138(n30138), .n23916(n23916), 
            .n25979(n25979), .clk_enable_222(clk_enable_222), .n26633(n26633), 
            .n30028(n30028), .n26779(n26779), .n30198(n30198), .n32(n32), 
            .\spi_data_r[1] (spi_data_r[1]), .\spi_data_r[2] (spi_data_r[2]), 
            .NSL(NSL), .EM_STOP(EM_STOP), .n25721(n25721), .n25547(n25547), 
            .n24169(n24169), .n18440(n18440), .n28402(n28402), .n28524(n28524), 
            .n30045(n30045), .n29999(n29999), .n28486(n28486), .\spi_addr_r[4] (spi_addr_r[4]), 
            .\spi_addr_r[2] (spi_addr_r[2]), .n27013(n27013), .\spi_cmd_r[0] (spi_cmd_r[0]), 
            .spi_data_valid_r(spi_data_valid_r), .\spi_addr_r[3] (spi_addr_r[3]), 
            .n30052(n30052), .n30007(n30007), .clk_enable_242(clk_enable_242), 
            .n29994(n29994), .n30199(n30199), .n25739(n25739), .n25699(n25699), 
            .n25941(n25941), .n25943(n25943), .n25801(n25801), .\spi_cmd_r[3] (spi_cmd_r[3]), 
            .n30044(n30044), .clk_enable_256(clk_enable_256), .\spi_cmd_r[1] (spi_cmd_r[1]), 
            .\spi_cmd_r[4] (spi_cmd_r[4]), .\spi_cmd_r[5] (spi_cmd_r[5]), 
            .reset_r(reset_r), .reset_r_N_4129(reset_r_N_4129), .n30043(n30043), 
            .mode_adj_653(mode_adj_7725), .n30018(n30018), .pin_io_out_4(pin_io_out_4), 
            .\pin_intrpt[2] (pin_intrpt[2]), .\quad_homing[0] (quad_homing[0]), 
            .n25869(n25869), .n30151(n30151)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(354[3] 397[2])
    \quad_decoder(DEV_ID=3)  \quad_ins_3..u_quad_decoder  (.n47(n47_adj_7734), 
            .clk(clk), .n30185(n30185), .\quad_b[3] (quad_b[3]), .\spi_data_out_r_39__N_1639[0] (spi_data_out_r_39__N_1639[0]), 
            .\pin_intrpt[11] (pin_intrpt[11]), .\quad_a[3] (quad_a[3]), 
            .quad_homing({quad_homing_adj_7853}), .clk_enable_687(clk_enable_687), 
            .\spi_data_r[0] (spi_data_r[0]), .clk_enable_727(clk_enable_727), 
            .spi_data_out_r_39__N_1679(spi_data_out_r_39__N_1679), .spi_data_out_r_39__N_1868(spi_data_out_r_39__N_1868), 
            .n29990(n29990), .\spi_data_out_r_39__N_1639[31] (spi_data_out_r_39__N_1639[31]), 
            .\spi_data_out_r_39__N_1639[30] (spi_data_out_r_39__N_1639[30]), 
            .\spi_data_out_r_39__N_1639[29] (spi_data_out_r_39__N_1639[29]), 
            .\spi_data_out_r_39__N_1639[28] (spi_data_out_r_39__N_1639[28]), 
            .\spi_data_out_r_39__N_1639[27] (spi_data_out_r_39__N_1639[27]), 
            .\spi_data_out_r_39__N_1639[26] (spi_data_out_r_39__N_1639[26]), 
            .\spi_data_out_r_39__N_1639[25] (spi_data_out_r_39__N_1639[25]), 
            .\spi_data_out_r_39__N_1639[24] (spi_data_out_r_39__N_1639[24]), 
            .\spi_data_out_r_39__N_1639[23] (spi_data_out_r_39__N_1639[23]), 
            .\spi_data_out_r_39__N_1639[22] (spi_data_out_r_39__N_1639[22]), 
            .\spi_data_out_r_39__N_1639[21] (spi_data_out_r_39__N_1639[21]), 
            .\spi_data_out_r_39__N_1639[20] (spi_data_out_r_39__N_1639[20]), 
            .\spi_data_out_r_39__N_1639[19] (spi_data_out_r_39__N_1639[19]), 
            .\spi_data_out_r_39__N_1639[18] (spi_data_out_r_39__N_1639[18]), 
            .\spi_data_out_r_39__N_1639[17] (spi_data_out_r_39__N_1639[17]), 
            .\spi_data_out_r_39__N_1639[16] (spi_data_out_r_39__N_1639[16]), 
            .\spi_data_out_r_39__N_1639[15] (spi_data_out_r_39__N_1639[15]), 
            .\spi_data_out_r_39__N_1639[14] (spi_data_out_r_39__N_1639[14]), 
            .\spi_data_out_r_39__N_1639[13] (spi_data_out_r_39__N_1639[13]), 
            .\spi_data_out_r_39__N_1639[12] (spi_data_out_r_39__N_1639[12]), 
            .\spi_data_out_r_39__N_1639[11] (spi_data_out_r_39__N_1639[11]), 
            .\spi_data_out_r_39__N_1639[10] (spi_data_out_r_39__N_1639[10]), 
            .\spi_data_out_r_39__N_1639[9] (spi_data_out_r_39__N_1639[9]), 
            .\spi_data_out_r_39__N_1639[8] (spi_data_out_r_39__N_1639[8]), 
            .\spi_data_out_r_39__N_1639[7] (spi_data_out_r_39__N_1639[7]), 
            .\spi_data_out_r_39__N_1639[6] (spi_data_out_r_39__N_1639[6]), 
            .\spi_data_out_r_39__N_1639[5] (spi_data_out_r_39__N_1639[5]), 
            .\spi_data_out_r_39__N_1639[4] (spi_data_out_r_39__N_1639[4]), 
            .\spi_data_out_r_39__N_1639[3] (spi_data_out_r_39__N_1639[3]), 
            .\spi_data_out_r_39__N_1639[2] (spi_data_out_r_39__N_1639[2]), 
            .\spi_data_out_r_39__N_1639[1] (spi_data_out_r_39__N_1639[1]), 
            .n1(n1_adj_7723), .\spi_data_r[1] (spi_data_r[1]), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[3] (spi_data_r[3]), .\spi_data_r[4] (spi_data_r[4]), 
            .\spi_data_r[5] (spi_data_r[5]), .\spi_data_r[6] (spi_data_r[6]), 
            .\spi_data_r[7] (spi_data_r[7]), .\spi_data_r[8] (spi_data_r[8]), 
            .\spi_data_r[9] (spi_data_r[9]), .\spi_data_r[10] (spi_data_r[10]), 
            .\spi_data_r[11] (spi_data_r[11]), .\spi_data_r[12] (spi_data_r[12]), 
            .\spi_data_r[13] (spi_data_r[13]), .\spi_data_r[14] (spi_data_r[14]), 
            .\spi_data_r[15] (spi_data_r[15]), .\spi_data_r[16] (spi_data_r[16]), 
            .\spi_data_r[17] (spi_data_r[17]), .\spi_data_r[18] (spi_data_r[18]), 
            .\spi_data_r[19] (spi_data_r[19]), .\spi_data_r[20] (spi_data_r[20]), 
            .\spi_data_r[21] (spi_data_r[21]), .\spi_data_r[22] (spi_data_r[22]), 
            .\spi_data_r[23] (spi_data_r[23]), .\spi_data_r[24] (spi_data_r[24]), 
            .\spi_data_r[25] (spi_data_r[25]), .\spi_data_r[26] (spi_data_r[26]), 
            .\spi_data_r[27] (spi_data_r[27]), .\spi_data_r[28] (spi_data_r[28]), 
            .\spi_data_r[29] (spi_data_r[29]), .\spi_data_r[30] (spi_data_r[30]), 
            .\spi_data_r[31] (spi_data_r[31]), .resetn_c(resetn_c), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(263[3] 283[2])
    \stepper(DEV_ID=3,UART_ADDRESS_WIDTH=4)  \stepper_ins_3..u_stepper  (.clk(clk), 
            .GND_net(GND_net), .reset_r(reset_r_adj_7679), .clk_enable_28(clk_enable_28), 
            .n30185(n30185), .n29995(n29995), .clk_1MHz(clk_1MHz), .clk_enable_178(clk_enable_178), 
            .\spi_data_r[0] (spi_data_r[0]), .n30188(n30188), .spi_data_out_r_39__N_4854({spi_data_out_r_39__N_4854}), 
            .\spi_data_out_r_39__N_5105[0] (spi_data_out_r_39__N_5105[0]), 
            .resetn_c(resetn_c), .\SLO_buf[0] (SLO_buf_adj_8193[0]), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[1] (spi_data_r[1]), .spi_data_out_r_39__N_4894(spi_data_out_r_39__N_4894), 
            .spi_data_out_r_39__N_5191(spi_data_out_r_39__N_5191), .digital_output_r(digital_output_r_adj_7680), 
            .clk_enable_254(clk_enable_254), .n28554(n28554), .pin_io_c_38(pin_io_c_38), 
            .\spi_data_out_r_39__N_5105[1] (spi_data_out_r_39__N_5105[1]), 
            .\spi_data_out_r_39__N_5105[2] (spi_data_out_r_39__N_5105[2]), 
            .\spi_data_out_r_39__N_5105[3] (spi_data_out_r_39__N_5105[3]), 
            .\spi_data_out_r_39__N_5105[4] (spi_data_out_r_39__N_5105[4]), 
            .\spi_data_out_r_39__N_5105[5] (spi_data_out_r_39__N_5105[5]), 
            .\spi_data_out_r_39__N_5105[6] (spi_data_out_r_39__N_5105[6]), 
            .\spi_data_out_r_39__N_5105[7] (spi_data_out_r_39__N_5105[7]), 
            .\spi_data_out_r_39__N_5105[8] (spi_data_out_r_39__N_5105[8]), 
            .\spi_data_out_r_39__N_5105[9] (spi_data_out_r_39__N_5105[9]), 
            .\spi_data_out_r_39__N_5105[10] (spi_data_out_r_39__N_5105[10]), 
            .\spi_data_out_r_39__N_5105[11] (spi_data_out_r_39__N_5105[11]), 
            .\spi_data_out_r_39__N_5105[12] (spi_data_out_r_39__N_5105[12]), 
            .\spi_data_out_r_39__N_5105[13] (spi_data_out_r_39__N_5105[13]), 
            .\spi_data_out_r_39__N_5105[14] (spi_data_out_r_39__N_5105[14]), 
            .\spi_data_out_r_39__N_5105[15] (spi_data_out_r_39__N_5105[15]), 
            .n29991(n29991), .\spi_data_out_r_39__N_5105[32] (spi_data_out_r_39__N_5105[32]), 
            .\spi_data_out_r_39__N_5105[33] (spi_data_out_r_39__N_5105[33]), 
            .\spi_data_out_r_39__N_5105[34] (spi_data_out_r_39__N_5105[34]), 
            .\spi_data_out_r_39__N_5105[35] (spi_data_out_r_39__N_5105[35]), 
            .\SLO_buf[10] (SLO_buf_adj_8193[10]), .\SLO_buf[11] (SLO_buf_adj_8193[11]), 
            .\SLO_buf[12] (SLO_buf_adj_8193[12]), .\SLO_buf[13] (SLO_buf_adj_8193[13]), 
            .\SLO_buf[1] (SLO_buf_adj_8193[1]), .\SLO_buf[2] (SLO_buf_adj_8193[2]), 
            .\SLO_buf[3] (SLO_buf_adj_8193[3]), .\SLO_buf[4] (SLO_buf_adj_8193[4]), 
            .\SLO_buf[5] (SLO_buf_adj_8193[5]), .\SLO_buf[6] (SLO_buf_adj_8193[6]), 
            .\SLO_buf[7] (SLO_buf_adj_8193[7]), .\SLO_buf[8] (SLO_buf_adj_8193[8]), 
            .\SLO_buf[9] (SLO_buf_adj_8193[9]), .\SLO_buf[14] (SLO_buf_adj_8193[14]), 
            .\SLO_buf[15] (SLO_buf_adj_8193[15]), .\SLO_buf[16] (SLO_buf_adj_8193[16]), 
            .\SLO_buf[17] (SLO_buf_adj_8193[17]), .\SLO_buf[18] (SLO_buf_adj_8193[18]), 
            .\SLO_buf[19] (SLO_buf_adj_8193[19]), .\SLO_buf[20] (SLO_buf_adj_8193[20]), 
            .\SLO_buf[21] (SLO_buf_adj_8193[21]), .\SLO_buf[22] (SLO_buf_adj_8193[22]), 
            .\SLO_buf[23] (SLO_buf_adj_8193[23]), .\SLO_buf[24] (SLO_buf_adj_8193[24]), 
            .\SLO_buf[25] (SLO_buf_adj_8193[25]), .\SLO_buf[26] (SLO_buf_adj_8193[26]), 
            .\SLO_buf[27] (SLO_buf_adj_8193[27]), .\SLO_buf[28] (SLO_buf_adj_8193[28]), 
            .\SLO_buf[29] (SLO_buf_adj_8193[29]), .NSL(NSL_adj_7681), .\quad_homing[0] (quad_homing_adj_7853[0]), 
            .pin_io_c_34(pin_io_c_34), .n25873(n25873), .mode(mode_adj_7728), 
            .\cs_decoded[6] (cs_decoded[6]), .n7170(n7170), .n30082(n30082), 
            .n7166(n7166), .n30091(n30091), .pin_io_out_35(pin_io_out_35), 
            .n29943(n29943), .pin_io_c_33(pin_io_c_33), .\pin_intrpt[10] (pin_intrpt[10]), 
            .pin_io_c_32(pin_io_c_32), .\pin_intrpt[9] (pin_intrpt[9]), 
            .\pin_intrpt[11] (pin_intrpt[11]), .n7269(n7269), .UC_TXD0_c(UC_TXD0_c), 
            .OW_ID_N_5147(OW_ID_N_5147), .n30050(n30050), .ENC_O_N_5155(ENC_O_N_5155), 
            .OW_ID_N_5153(OW_ID_N_5153), .\quad_a[3] (quad_a[3]), .pin_io_out_39(pin_io_out_39), 
            .\quad_b[3] (quad_b[3]), .\uart_slot_en[1] (uart_slot_en[1]), 
            .\uart_slot_en[0] (uart_slot_en[0]), .n10696(n10696), .mode_adj_652(mode_adj_7729), 
            .tx_N_6586(tx_N_6586)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(354[3] 397[2])
    \stepper(DEV_ID=4,UART_ADDRESS_WIDTH=4)  \stepper_ins_4..u_stepper  (.reset_r(reset_r_adj_7713), 
            .clk(clk), .n30185(n30185), .n30031(n30031), .clk_1MHz(clk_1MHz), 
            .GND_net(GND_net), .n30146(n30146), .clk_enable_641(clk_enable_641), 
            .\spi_data_r[0] (spi_data_r[0]), .spi_data_out_r_39__N_5197({spi_data_out_r_39__N_5197}), 
            .resetn_c(resetn_c), .digital_output_r(digital_output_r_adj_7714), 
            .n28549(n28549), .\uart_slot_en[0] (uart_slot_en[0]), .n30091(n30091), 
            .n29594(n29594), .spi_data_out_r_39__N_5237(spi_data_out_r_39__N_5237), 
            .spi_data_out_r_39__N_5534(spi_data_out_r_39__N_5534), .pin_io_out_45(pin_io_out_45), 
            .\uart_slot_en[2] (uart_slot_en[2]), .n29481(n29481), .pin_io_c_48(pin_io_c_48), 
            .\spi_data_r[1] (spi_data_r[1]), .\spi_data_r[2] (spi_data_r[2]), 
            .n47(n47), .NSL(NSL_adj_7715), .n25979(n25979), .n23916(n23916), 
            .n30199(n30199), .\quad_homing[0] (quad_homing_adj_7891[0]), 
            .pin_io_c_44(pin_io_c_44), .n25893(n25893), .ENC_O_N_5498(ENC_O_N_5498), 
            .n30180(n30180), .TX_IN_N_6565(TX_IN_N_6565), .n7163(n7163), 
            .\uart_slot_en[1] (uart_slot_en[1]), .n23722(n23722), .EM_STOP(EM_STOP), 
            .n25699(n25699), .UC_TXD0_c(UC_TXD0_c), .OW_ID_N_5490(OW_ID_N_5490), 
            .n30050(n30050), .n30120(n30120), .pin_io_out_49(pin_io_out_49), 
            .\quad_b[4] (quad_b[4]), .\quad_a[4] (quad_a[4]), .\pin_intrpt[14] (pin_intrpt[14]), 
            .n30055(n30055), .OW_ID_N_5496(OW_ID_N_5496), .n7266(n7266), 
            .pin_io_c_42(pin_io_c_42), .\pin_intrpt[12] (pin_intrpt[12]), 
            .pin_io_c_43(pin_io_c_43), .\pin_intrpt[13] (pin_intrpt[13])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(354[3] 397[2])
    spi_slave_top spi_slave_top_inst (.spi_addr_r({spi_addr_r}), .clk(clk), 
            .n30080(n30080), .n30185(n30185), .spi_data_valid_r(spi_data_valid_r), 
            .spi_data_valid(spi_data_valid), .n23916(n23916), .n30035(n30035), 
            .\spi_data_r[0] (spi_data_r[0]), .clk_enable_161(clk_enable_161), 
            .spi_scsn_c(spi_scsn_c), .spi_addr_valid(spi_addr_valid), .spi_cmd_valid(spi_cmd_valid), 
            .\spi_data_r[31] (spi_data_r[31]), .\spi_data_r[30] (spi_data_r[30]), 
            .\spi_data_r[29] (spi_data_r[29]), .\spi_data_r[28] (spi_data_r[28]), 
            .\spi_data_r[27] (spi_data_r[27]), .\spi_data_r[26] (spi_data_r[26]), 
            .\spi_data_r[25] (spi_data_r[25]), .\spi_data_r[24] (spi_data_r[24]), 
            .\spi_data_r[23] (spi_data_r[23]), .\spi_data_r[22] (spi_data_r[22]), 
            .\spi_data_r[21] (spi_data_r[21]), .\spi_data_r[20] (spi_data_r[20]), 
            .\spi_data_r[19] (spi_data_r[19]), .\spi_data_r[18] (spi_data_r[18]), 
            .\spi_data_r[17] (spi_data_r[17]), .\spi_data_r[16] (spi_data_r[16]), 
            .spi_cmd_r({spi_cmd_r}), .n28328(n28328), .n26327(n26327), 
            .\spi_data_r[15] (spi_data_r[15]), .\spi_data_r[14] (spi_data_r[14]), 
            .\spi_data_r[13] (spi_data_r[13]), .\spi_data_r[12] (spi_data_r[12]), 
            .\spi_data_r[11] (spi_data_r[11]), .\spi_data_r[10] (spi_data_r[10]), 
            .\spi_data_r[9] (spi_data_r[9]), .\spi_data_r[8] (spi_data_r[8]), 
            .\spi_data_r[7] (spi_data_r[7]), .\spi_data_r[6] (spi_data_r[6]), 
            .\spi_data_r[5] (spi_data_r[5]), .\spi_data_r[4] (spi_data_r[4]), 
            .\spi_data_r[3] (spi_data_r[3]), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[1] (spi_data_r[1]), .\spi_data_out_r[0] (spi_data_out_r[0]), 
            .n26621(n26621), .n26819(n26819), .n27013(n27013), .n27015(n27015), 
            .n30144(n30144), .n30155(n30155), .n18440(n18440), .n28524(n28524), 
            .n4(n4_adj_7388), .n30044(n30044), .n23526(n23526), .n26545(n26545), 
            .n30151(n30151), .n30094(n30094), .quad_set_valid_N_1158(quad_set_valid_N_1158), 
            .n23732(n23732), .n26497(n26497), .n30209(n30209), .n28260(n28260), 
            .n30214(n30214), .\spi_cmd[2] (spi_cmd[2]), .\spi_data_out_r[1] (spi_data_out_r[1]), 
            .\spi_data_out_r[3] (spi_data_out_r[3]), .\spi_data_out_r[4] (spi_data_out_r[4]), 
            .\spi_data_out_r[5] (spi_data_out_r[5]), .\spi_data_out_r[6] (spi_data_out_r[6]), 
            .\spi_data_out_r[7] (spi_data_out_r[7]), .\spi_data_out_r_39__N_5197[8] (spi_data_out_r_39__N_5197[8]), 
            .n16(n16_adj_7461), .spi_data_out_r_39__N_5237(spi_data_out_r_39__N_5237), 
            .\spi_data_out_r[10] (spi_data_out_r[10]), .\spi_data_out_r[11] (spi_data_out_r[11]), 
            .\spi_data_out_r[12] (spi_data_out_r[12]), .\spi_data_out_r[13] (spi_data_out_r[13]), 
            .\spi_data_out_r[14] (spi_data_out_r[14]), .\spi_data_out_r[15] (spi_data_out_r[15]), 
            .\spi_data_out_r[16] (spi_data_out_r[16]), .\spi_data_out_r[17] (spi_data_out_r[17]), 
            .\spi_data_out_r[18] (spi_data_out_r[18]), .\spi_data_out_r[19] (spi_data_out_r[19]), 
            .\spi_data_out_r[20] (spi_data_out_r[20]), .\spi_data_out_r[21] (spi_data_out_r[21]), 
            .\spi_data_out_r[22] (spi_data_out_r[22]), .\spi_data_out_r[23] (spi_data_out_r[23]), 
            .\spi_data_out_r[24] (spi_data_out_r[24]), .\spi_data_out_r[25] (spi_data_out_r[25]), 
            .\spi_data_out_r[26] (spi_data_out_r[26]), .\spi_data_out_r[27] (spi_data_out_r[27]), 
            .\spi_data_out_r[28] (spi_data_out_r[28]), .\spi_data_out_r[29] (spi_data_out_r[29]), 
            .\spi_data_out_r[30] (spi_data_out_r[30]), .\spi_data_out_r[31] (spi_data_out_r[31]), 
            .\spi_data_out_r[32] (spi_data_out_r[32]), .\spi_data_out_r[33] (spi_data_out_r[33]), 
            .\spi_data_out_r[34] (spi_data_out_r[34]), .\spi_data_out_r[35] (spi_data_out_r[35]), 
            .\spi_data_out_r[36] (spi_data_out_r[36]), .\spi_data_out_r[37] (spi_data_out_r[37]), 
            .\spi_data_out_r[38] (spi_data_out_r[38]), .\spi_data_out_r[39] (spi_data_out_r[39]), 
            .\spi_data_out_r_39__N_5540[8] (spi_data_out_r_39__N_5540[8]), 
            .n18(n18_adj_7460), .spi_data_out_r_39__N_5580(spi_data_out_r_39__N_5580), 
            .\spi_data_out_r_39__N_4168[8] (spi_data_out_r_39__N_4168[8]), 
            .n3(n3), .spi_data_out_r_39__N_4208(spi_data_out_r_39__N_4208), 
            .\spi_data_out_r_39__N_5883[8] (spi_data_out_r_39__N_5883[8]), 
            .\spi_data_out_r_39__N_4854[8] (spi_data_out_r_39__N_4854[8]), 
            .spi_data_out_r_39__N_5923(spi_data_out_r_39__N_5923), .spi_data_out_r_39__N_4894(spi_data_out_r_39__N_4894), 
            .\spi_data_out_r_39__N_2109[8] (spi_data_out_r_39__N_2109[8]), 
            .n5(n5_adj_7462), .spi_data_out_r_39__N_2149(spi_data_out_r_39__N_2149), 
            .\spi_data_out_r_39__N_1404[8] (spi_data_out_r_39__N_1404[8]), 
            .\spi_data_out_r_39__N_934[8] (spi_data_out_r_39__N_934[8]), .spi_data_out_r_39__N_1444(spi_data_out_r_39__N_1444), 
            .spi_data_out_r_39__N_974(spi_data_out_r_39__N_974), .n28384(n28384), 
            .\spi_data_out_r_39__N_2344[8] (spi_data_out_r_39__N_2344[8]), 
            .\spi_data_out_r_39__N_1874[8] (spi_data_out_r_39__N_1874[8]), 
            .spi_data_out_r_39__N_2384(spi_data_out_r_39__N_2384), .spi_data_out_r_39__N_1914(spi_data_out_r_39__N_1914), 
            .\spi_data_out_r_39__N_4168[9] (spi_data_out_r_39__N_4168[9]), 
            .n16_adj_329(n16), .\spi_data_out_r_39__N_5883[9] (spi_data_out_r_39__N_5883[9]), 
            .n21(n21), .\spi_data_out_r_39__N_4854[9] (spi_data_out_r_39__N_4854[9]), 
            .n2(n2), .\spi_data_out_r_39__N_5197[9] (spi_data_out_r_39__N_5197[9]), 
            .\spi_data_out_r_39__N_4511[9] (spi_data_out_r_39__N_4511[9]), 
            .spi_data_out_r_39__N_4551(spi_data_out_r_39__N_4551), .\spi_data_out_r_39__N_1874[9] (spi_data_out_r_39__N_1874[9]), 
            .n5_adj_330(n5), .\spi_data_out_r_39__N_2344[9] (spi_data_out_r_39__N_2344[9]), 
            .\spi_data_out_r_39__N_2109[9] (spi_data_out_r_39__N_2109[9]), 
            .\spi_data_out_r_39__N_1404[9] (spi_data_out_r_39__N_1404[9]), 
            .\spi_data_out_r_39__N_1169[9] (spi_data_out_r_39__N_1169[9]), 
            .spi_data_out_r_39__N_1209(spi_data_out_r_39__N_1209), .n21_adj_331(n21_adj_7670), 
            .n19(n19), .\spi_data_out_r_39__N_5197[2] (spi_data_out_r_39__N_5197[2]), 
            .n22(n22), .\spi_data_out_r_39__N_2863[2] (spi_data_out_r_39__N_2863[2]), 
            .\spi_data_out_r_39__N_2721[2] (spi_data_out_r_39__N_2721[2]), 
            .clear_intrpt(clear_intrpt_adj_7664), .clear_intrpt_adj_332(clear_intrpt_adj_7662), 
            .\spi_data_out_r_39__N_4511[2] (spi_data_out_r_39__N_4511[2]), 
            .\spi_data_out_r_39__N_4168[2] (spi_data_out_r_39__N_4168[2]), 
            .\spi_data_out_r_39__N_3005[2] (spi_data_out_r_39__N_3005[2]), 
            .n14(n14), .n9(n9), .clear_intrpt_adj_333(clear_intrpt_adj_7666), 
            .\spi_data_out_r_39__N_2792[2] (spi_data_out_r_39__N_2792[2]), 
            .\spi_data_out_r_39__N_2650[2] (spi_data_out_r_39__N_2650[2]), 
            .clear_intrpt_adj_334(clear_intrpt_adj_7663), .clear_intrpt_adj_335(clear_intrpt_adj_7661), 
            .\spi_data_out_r_39__N_1169[2] (spi_data_out_r_39__N_1169[2]), 
            .n7(n7), .\spi_data_out_r_39__N_1639[2] (spi_data_out_r_39__N_1639[2]), 
            .\spi_data_out_r_39__N_1404[2] (spi_data_out_r_39__N_1404[2]), 
            .spi_data_out_r_39__N_1679(spi_data_out_r_39__N_1679), .\spi_data_out_r_39__N_1874[2] (spi_data_out_r_39__N_1874[2]), 
            .\spi_data_out_r_39__N_2344[2] (spi_data_out_r_39__N_2344[2]), 
            .\spi_data_out_r_39__N_3825[2] (spi_data_out_r_39__N_3825[2]), 
            .\spi_data_out_r_39__N_934[2] (spi_data_out_r_39__N_934[2]), .spi_data_out_r_39__N_3865(spi_data_out_r_39__N_3865), 
            .n25721(n25721), .n28358(n28358), .n26435(n26435), .n26521(n26521), 
            .n30090(n30090), .n26569(n26569), .n24066(n24066), .n28340(n28340), 
            .quad_set_valid_N_1393(quad_set_valid_N_1393), .n30071(n30071), 
            .n25571(n25571), .n26243(n26243), .n30062(n30062), .n25859(n25859), 
            .resetn_c(resetn_c), .n30210(n30210), .n30213(n30213), .n30023(n30023), 
            .n29995(n29995), .n29996(n29996), .clk_enable_254(clk_enable_254), 
            .clk_enable_259(clk_enable_259), .n30070(n30070), .n29993(n29993), 
            .n25643(n25643), .n30064(n30064), .n23537(n23537), .n31069(n31069), 
            .GND_net(GND_net), .spi_mosi_oe(spi_mosi_oe), .spi_mosi_o(spi_mosi_o), 
            .spi_miso_oe(spi_miso_oe), .spi_miso_o(spi_miso_o), .spi_clk_oe(spi_clk_oe), 
            .spi_clk_o(spi_clk_o), .spi_mosi_i(spi_mosi_i), .spi_miso_i(spi_miso_i), 
            .spi_clk_i(spi_clk_i), .VCC_net(VCC_net), .quad_buffer({quad_buffer}), 
            .quad_count({quad_count}), .\spi_data_out_r_39__N_1083[31] (spi_data_out_r_39__N_1083[31]), 
            .\spi_data_out_r_39__N_1083[29] (spi_data_out_r_39__N_1083[29]), 
            .\spi_data_out_r_39__N_1083[19] (spi_data_out_r_39__N_1083[19]), 
            .\spi_data_out_r_39__N_1083[18] (spi_data_out_r_39__N_1083[18]), 
            .quad_buffer_adj_644({quad_buffer_adj_7893}), .quad_count_adj_645({quad_count_adj_7892}), 
            .\spi_data_out_r_39__N_2023[26] (spi_data_out_r_39__N_2023[26]), 
            .n30198(n30198), .n32(n32), .clear_intrpt_N_2717(clear_intrpt_N_2717), 
            .n47(n47_adj_7732), .clear_intrpt_N_2930(clear_intrpt_N_2930), 
            .clear_intrpt_N_2788(clear_intrpt_N_2788), .clear_intrpt_N_2859(clear_intrpt_N_2859), 
            .n47_adj_400(n47_adj_7731), .quad_buffer_adj_646({quad_buffer_adj_7969}), 
            .quad_count_adj_647({quad_count_adj_7968}), .\spi_data_out_r_39__N_2493[29] (spi_data_out_r_39__N_2493[29]), 
            .\spi_data_out_r_39__N_2493[28] (spi_data_out_r_39__N_2493[28]), 
            .\spi_data_out_r_39__N_2493[27] (spi_data_out_r_39__N_2493[27]), 
            .\spi_data_out_r_39__N_2493[26] (spi_data_out_r_39__N_2493[26]), 
            .n29997(n29997), .n29991(n29991), .\spi_data_out_r_39__N_2493[25] (spi_data_out_r_39__N_2493[25]), 
            .\spi_data_out_r_39__N_2493[24] (spi_data_out_r_39__N_2493[24]), 
            .\spi_data_out_r_39__N_2493[23] (spi_data_out_r_39__N_2493[23]), 
            .\spi_data_out_r_39__N_2493[22] (spi_data_out_r_39__N_2493[22]), 
            .\spi_data_out_r_39__N_2493[21] (spi_data_out_r_39__N_2493[21]), 
            .\spi_data_out_r_39__N_2493[20] (spi_data_out_r_39__N_2493[20]), 
            .\spi_data_out_r_39__N_2493[19] (spi_data_out_r_39__N_2493[19]), 
            .\spi_data_out_r_39__N_2493[18] (spi_data_out_r_39__N_2493[18]), 
            .\spi_data_out_r_39__N_2493[17] (spi_data_out_r_39__N_2493[17]), 
            .\spi_data_out_r_39__N_2493[16] (spi_data_out_r_39__N_2493[16]), 
            .\spi_data_out_r_39__N_2493[15] (spi_data_out_r_39__N_2493[15]), 
            .\spi_data_out_r_39__N_2493[14] (spi_data_out_r_39__N_2493[14]), 
            .\spi_data_out_r_39__N_2493[13] (spi_data_out_r_39__N_2493[13]), 
            .\spi_data_out_r_39__N_2493[12] (spi_data_out_r_39__N_2493[12]), 
            .\spi_data_out_r_39__N_2493[11] (spi_data_out_r_39__N_2493[11]), 
            .\spi_data_out_r_39__N_2493[10] (spi_data_out_r_39__N_2493[10]), 
            .\spi_data_out_r_39__N_2493[9] (spi_data_out_r_39__N_2493[9]), 
            .\spi_data_out_r_39__N_2493[8] (spi_data_out_r_39__N_2493[8]), 
            .\spi_data_out_r_39__N_2493[7] (spi_data_out_r_39__N_2493[7]), 
            .\spi_data_out_r_39__N_1083[9] (spi_data_out_r_39__N_1083[9]), 
            .\spi_data_out_r_39__N_1083[8] (spi_data_out_r_39__N_1083[8]), 
            .\spi_data_out_r_39__N_2493[6] (spi_data_out_r_39__N_2493[6]), 
            .\spi_data_out_r_39__N_2493[5] (spi_data_out_r_39__N_2493[5]), 
            .\spi_data_out_r_39__N_2493[4] (spi_data_out_r_39__N_2493[4]), 
            .\spi_data_out_r_39__N_2493[3] (spi_data_out_r_39__N_2493[3]), 
            .\spi_data_out_r_39__N_2493[2] (spi_data_out_r_39__N_2493[2]), 
            .\spi_data_out_r_39__N_2493[1] (spi_data_out_r_39__N_2493[1]), 
            .\spi_data_out_r_39__N_2023[20] (spi_data_out_r_39__N_2023[20]), 
            .quad_buffer_adj_648({quad_buffer_adj_7931}), .quad_count_adj_649({quad_count_adj_7930}), 
            .\spi_data_out_r_39__N_2258[0] (spi_data_out_r_39__N_2258[0]), 
            .\spi_data_out_r_39__N_2258[31] (spi_data_out_r_39__N_2258[31]), 
            .\spi_data_out_r_39__N_2258[30] (spi_data_out_r_39__N_2258[30]), 
            .\spi_data_out_r_39__N_2258[29] (spi_data_out_r_39__N_2258[29]), 
            .\spi_data_out_r_39__N_2258[28] (spi_data_out_r_39__N_2258[28]), 
            .\spi_data_out_r_39__N_2258[27] (spi_data_out_r_39__N_2258[27]), 
            .\spi_data_out_r_39__N_2258[26] (spi_data_out_r_39__N_2258[26]), 
            .n26779(n26779), .\spi_data_out_r_39__N_2258[25] (spi_data_out_r_39__N_2258[25]), 
            .\spi_data_out_r_39__N_2258[24] (spi_data_out_r_39__N_2258[24]), 
            .\spi_data_out_r_39__N_1083[22] (spi_data_out_r_39__N_1083[22]), 
            .\spi_data_out_r_39__N_2258[23] (spi_data_out_r_39__N_2258[23]), 
            .\spi_data_out_r_39__N_2258[22] (spi_data_out_r_39__N_2258[22]), 
            .\spi_data_out_r_39__N_2258[21] (spi_data_out_r_39__N_2258[21]), 
            .\spi_data_out_r_39__N_2258[20] (spi_data_out_r_39__N_2258[20]), 
            .\spi_data_out_r_39__N_2258[19] (spi_data_out_r_39__N_2258[19]), 
            .\spi_data_out_r_39__N_2258[18] (spi_data_out_r_39__N_2258[18]), 
            .n47_adj_529(n47), .\spi_data_out_r_39__N_2258[17] (spi_data_out_r_39__N_2258[17]), 
            .\spi_data_out_r_39__N_2258[16] (spi_data_out_r_39__N_2258[16]), 
            .\spi_data_out_r_39__N_2258[15] (spi_data_out_r_39__N_2258[15]), 
            .\spi_data_out_r_39__N_2258[14] (spi_data_out_r_39__N_2258[14]), 
            .\spi_data_out_r_39__N_2258[13] (spi_data_out_r_39__N_2258[13]), 
            .\spi_data_out_r_39__N_2258[12] (spi_data_out_r_39__N_2258[12]), 
            .\spi_data_out_r_39__N_2258[11] (spi_data_out_r_39__N_2258[11]), 
            .\spi_data_out_r_39__N_2258[10] (spi_data_out_r_39__N_2258[10]), 
            .\spi_data_out_r_39__N_2258[9] (spi_data_out_r_39__N_2258[9]), 
            .n30019(n30019), .n47_adj_530(n47_adj_7716), .\spi_data_out_r_39__N_2258[8] (spi_data_out_r_39__N_2258[8]), 
            .\spi_data_out_r_39__N_2258[7] (spi_data_out_r_39__N_2258[7]), 
            .n30027(n30027), .n47_adj_531(n47_adj_7730), .\spi_data_out_r_39__N_2258[6] (spi_data_out_r_39__N_2258[6]), 
            .\spi_data_out_r_39__N_2258[5] (spi_data_out_r_39__N_2258[5]), 
            .\spi_data_out_r_39__N_2258[4] (spi_data_out_r_39__N_2258[4]), 
            .\spi_data_out_r_39__N_2258[3] (spi_data_out_r_39__N_2258[3]), 
            .\spi_data_out_r_39__N_1083[17] (spi_data_out_r_39__N_1083[17]), 
            .\spi_data_out_r_39__N_2258[2] (spi_data_out_r_39__N_2258[2]), 
            .\spi_data_out_r_39__N_2023[19] (spi_data_out_r_39__N_2023[19]), 
            .\spi_data_out_r_39__N_2258[1] (spi_data_out_r_39__N_2258[1]), 
            .\SLO_buf[4] (SLO_buf_adj_8193[4]), .\SLO_buf[14] (SLO_buf_adj_8193[14]), 
            .\spi_data_out_r_39__N_5105[0] (spi_data_out_r_39__N_5105[0]), 
            .\SLO_buf[3] (SLO_buf_adj_8193[3]), .\SLO_buf[9] (SLO_buf_adj_8193[9]), 
            .\spi_data_out_r_39__N_5105[35] (spi_data_out_r_39__N_5105[35]), 
            .\SLO_buf[2] (SLO_buf_adj_8193[2]), .\SLO_buf[8] (SLO_buf_adj_8193[8]), 
            .\spi_data_out_r_39__N_5105[34] (spi_data_out_r_39__N_5105[34]), 
            .\SLO_buf[1] (SLO_buf_adj_8193[1]), .\SLO_buf[7] (SLO_buf_adj_8193[7]), 
            .\spi_data_out_r_39__N_5105[33] (spi_data_out_r_39__N_5105[33]), 
            .quad_buffer_adj_650({quad_buffer_adj_7817}), .quad_count_adj_651({quad_count_adj_7816}), 
            .\spi_data_out_r_39__N_1553[0] (spi_data_out_r_39__N_1553[0]), 
            .\spi_data_out_r_39__N_1553[31] (spi_data_out_r_39__N_1553[31]), 
            .\SLO_buf[0] (SLO_buf_adj_8193[0]), .\SLO_buf[6] (SLO_buf_adj_8193[6]), 
            .\spi_data_out_r_39__N_5105[32] (spi_data_out_r_39__N_5105[32]), 
            .\SLO_buf[19] (SLO_buf_adj_8193[19]), .\SLO_buf[29] (SLO_buf_adj_8193[29]), 
            .\spi_data_out_r_39__N_5105[15] (spi_data_out_r_39__N_5105[15]), 
            .\spi_data_out_r_39__N_1553[30] (spi_data_out_r_39__N_1553[30]), 
            .\spi_data_out_r_39__N_1553[29] (spi_data_out_r_39__N_1553[29]), 
            .\spi_data_out_r_39__N_1553[28] (spi_data_out_r_39__N_1553[28]), 
            .\spi_data_out_r_39__N_1553[27] (spi_data_out_r_39__N_1553[27]), 
            .\SLO_buf[18] (SLO_buf_adj_8193[18]), .\SLO_buf[28] (SLO_buf_adj_8193[28]), 
            .\spi_data_out_r_39__N_5105[14] (spi_data_out_r_39__N_5105[14]), 
            .\spi_data_out_r_39__N_1553[26] (spi_data_out_r_39__N_1553[26]), 
            .\SLO_buf[17] (SLO_buf_adj_8193[17]), .\SLO_buf[27] (SLO_buf_adj_8193[27]), 
            .\spi_data_out_r_39__N_5105[13] (spi_data_out_r_39__N_5105[13]), 
            .\spi_data_out_r_39__N_2023[25] (spi_data_out_r_39__N_2023[25]), 
            .\spi_data_out_r_39__N_1553[25] (spi_data_out_r_39__N_1553[25]), 
            .\spi_data_out_r_39__N_1553[24] (spi_data_out_r_39__N_1553[24]), 
            .\SLO_buf[16] (SLO_buf_adj_8193[16]), .\SLO_buf[26] (SLO_buf_adj_8193[26]), 
            .\spi_data_out_r_39__N_5105[12] (spi_data_out_r_39__N_5105[12]), 
            .\spi_data_out_r_39__N_1553[23] (spi_data_out_r_39__N_1553[23]), 
            .\SLO_buf[15] (SLO_buf_adj_8193[15]), .\SLO_buf[25] (SLO_buf_adj_8193[25]), 
            .\spi_data_out_r_39__N_5105[11] (spi_data_out_r_39__N_5105[11]), 
            .\SLO_buf[24] (SLO_buf_adj_8193[24]), .\spi_data_out_r_39__N_5105[10] (spi_data_out_r_39__N_5105[10]), 
            .\spi_data_out_r_39__N_1553[22] (spi_data_out_r_39__N_1553[22]), 
            .\SLO_buf[13] (SLO_buf_adj_8193[13]), .\SLO_buf[23] (SLO_buf_adj_8193[23]), 
            .\spi_data_out_r_39__N_5105[9] (spi_data_out_r_39__N_5105[9]), 
            .\spi_data_out_r_39__N_1553[21] (spi_data_out_r_39__N_1553[21]), 
            .\spi_data_out_r_39__N_1553[20] (spi_data_out_r_39__N_1553[20]), 
            .\spi_data_out_r_39__N_1553[19] (spi_data_out_r_39__N_1553[19]), 
            .\spi_data_out_r_39__N_1553[18] (spi_data_out_r_39__N_1553[18]), 
            .\spi_data_out_r_39__N_1553[17] (spi_data_out_r_39__N_1553[17]), 
            .\spi_data_out_r_39__N_1553[16] (spi_data_out_r_39__N_1553[16]), 
            .\spi_data_out_r_39__N_1083[16] (spi_data_out_r_39__N_1083[16]), 
            .\spi_data_out_r_39__N_1553[15] (spi_data_out_r_39__N_1553[15]), 
            .\spi_data_out_r_39__N_1553[14] (spi_data_out_r_39__N_1553[14]), 
            .\spi_data_out_r_39__N_1553[13] (spi_data_out_r_39__N_1553[13]), 
            .\spi_data_out_r_39__N_1083[15] (spi_data_out_r_39__N_1083[15]), 
            .\SLO_buf[12] (SLO_buf_adj_8193[12]), .\SLO_buf[22] (SLO_buf_adj_8193[22]), 
            .\spi_data_out_r_39__N_5105[8] (spi_data_out_r_39__N_5105[8]), 
            .\spi_data_out_r_39__N_1553[12] (spi_data_out_r_39__N_1553[12]), 
            .\SLO_buf[11] (SLO_buf_adj_8193[11]), .\SLO_buf[21] (SLO_buf_adj_8193[21]), 
            .\spi_data_out_r_39__N_5105[7] (spi_data_out_r_39__N_5105[7]), 
            .\spi_data_out_r_39__N_1553[11] (spi_data_out_r_39__N_1553[11]), 
            .\SLO_buf[10] (SLO_buf_adj_8193[10]), .\SLO_buf[20] (SLO_buf_adj_8193[20]), 
            .\spi_data_out_r_39__N_5105[6] (spi_data_out_r_39__N_5105[6]), 
            .\spi_data_out_r_39__N_5105[5] (spi_data_out_r_39__N_5105[5]), 
            .\spi_data_out_r_39__N_1553[10] (spi_data_out_r_39__N_1553[10]), 
            .\spi_data_out_r_39__N_5105[4] (spi_data_out_r_39__N_5105[4]), 
            .\spi_data_out_r_39__N_1553[9] (spi_data_out_r_39__N_1553[9]), 
            .\spi_data_out_r_39__N_1553[8] (spi_data_out_r_39__N_1553[8]), 
            .\spi_data_out_r_39__N_1553[7] (spi_data_out_r_39__N_1553[7]), 
            .\spi_data_out_r_39__N_1553[6] (spi_data_out_r_39__N_1553[6]), 
            .\spi_data_out_r_39__N_5105[3] (spi_data_out_r_39__N_5105[3]), 
            .\spi_data_out_r_39__N_1553[5] (spi_data_out_r_39__N_1553[5]), 
            .\spi_data_out_r_39__N_1553[4] (spi_data_out_r_39__N_1553[4]), 
            .\spi_data_out_r_39__N_1553[3] (spi_data_out_r_39__N_1553[3]), 
            .\spi_data_out_r_39__N_2023[18] (spi_data_out_r_39__N_2023[18]), 
            .\spi_data_out_r_39__N_1553[2] (spi_data_out_r_39__N_1553[2]), 
            .\spi_data_out_r_39__N_1553[1] (spi_data_out_r_39__N_1553[1]), 
            .n47_adj_596(n47_adj_7735), .\spi_data_out_r_39__N_5105[2] (spi_data_out_r_39__N_5105[2]), 
            .\SLO_buf[5] (SLO_buf_adj_8193[5]), .\spi_data_out_r_39__N_5105[1] (spi_data_out_r_39__N_5105[1]), 
            .spi_data_out_r_39__N_2338(spi_data_out_r_39__N_2338), .n47_adj_597(n47_adj_7734), 
            .\spi_data_out_r_39__N_1083[14] (spi_data_out_r_39__N_1083[14]), 
            .\spi_data_out_r_39__N_1083[13] (spi_data_out_r_39__N_1083[13]), 
            .n30102(n30102), .\SLO_buf[4]_adj_598 (SLO_buf_adj_8127[4]), 
            .\SLO_buf[14]_adj_599 (SLO_buf_adj_8127[14]), .\spi_data_out_r_39__N_4419[0] (spi_data_out_r_39__N_4419[0]), 
            .\SLO_buf[3]_adj_600 (SLO_buf_adj_8127[3]), .\SLO_buf[9]_adj_601 (SLO_buf_adj_8127[9]), 
            .\spi_data_out_r_39__N_4419[35] (spi_data_out_r_39__N_4419[35]), 
            .spi_data_out_r_39__N_4505(spi_data_out_r_39__N_4505), .\spi_data_out_r_39__N_2023[17] (spi_data_out_r_39__N_2023[17]), 
            .\spi_data_out_r_39__N_2023[16] (spi_data_out_r_39__N_2023[16]), 
            .\spi_data_out_r_39__N_1083[7] (spi_data_out_r_39__N_1083[7]), 
            .\spi_data_out_r_39__N_1083[6] (spi_data_out_r_39__N_1083[6]), 
            .\spi_data_out_r_39__N_1083[20] (spi_data_out_r_39__N_1083[20]), 
            .\spi_data_out_r_39__N_2023[15] (spi_data_out_r_39__N_2023[15]), 
            .\status_cntr[12] (status_cntr[12]), .n25212(n25212), .\SLO_buf[2]_adj_602 (SLO_buf_adj_8127[2]), 
            .\SLO_buf[8]_adj_603 (SLO_buf_adj_8127[8]), .\spi_data_out_r_39__N_4419[34] (spi_data_out_r_39__N_4419[34]), 
            .\spi_data_out_r_39__N_2023[14] (spi_data_out_r_39__N_2023[14]), 
            .\SLO_buf[1]_adj_604 (SLO_buf_adj_8127[1]), .\SLO_buf[7]_adj_605 (SLO_buf_adj_8127[7]), 
            .\spi_data_out_r_39__N_4419[33] (spi_data_out_r_39__N_4419[33]), 
            .\SLO_buf[0]_adj_606 (SLO_buf_adj_8127[0]), .\SLO_buf[6]_adj_607 (SLO_buf_adj_8127[6]), 
            .\spi_data_out_r_39__N_4419[32] (spi_data_out_r_39__N_4419[32]), 
            .clear_intrpt_N_3072(clear_intrpt_N_3072), .\spi_data_out_r_39__N_2023[13] (spi_data_out_r_39__N_2023[13]), 
            .\SLO_buf[19]_adj_608 (SLO_buf_adj_8127[19]), .\SLO_buf[29]_adj_609 (SLO_buf_adj_8127[29]), 
            .\spi_data_out_r_39__N_4419[15] (spi_data_out_r_39__N_4419[15]), 
            .\spi_data_out_r_39__N_1083[5] (spi_data_out_r_39__N_1083[5]), 
            .\spi_data_out_r_39__N_1083[4] (spi_data_out_r_39__N_1083[4]), 
            .\spi_data_out_r_39__N_2023[12] (spi_data_out_r_39__N_2023[12]), 
            .\SLO_buf[18]_adj_610 (SLO_buf_adj_8127[18]), .\SLO_buf[28]_adj_611 (SLO_buf_adj_8127[28]), 
            .\spi_data_out_r_39__N_4419[14] (spi_data_out_r_39__N_4419[14]), 
            .\SLO_buf[17]_adj_612 (SLO_buf_adj_8127[17]), .\SLO_buf[27]_adj_613 (SLO_buf_adj_8127[27]), 
            .\spi_data_out_r_39__N_4419[13] (spi_data_out_r_39__N_4419[13]), 
            .\spi_data_out_r_39__N_1083[12] (spi_data_out_r_39__N_1083[12]), 
            .spi_data_out_r_39__N_4848(spi_data_out_r_39__N_4848), .\spi_data_out_r_39__N_1083[3] (spi_data_out_r_39__N_1083[3]), 
            .\spi_data_out_r_39__N_1083[2] (spi_data_out_r_39__N_1083[2]), 
            .\spi_data_out_r_39__N_2023[11] (spi_data_out_r_39__N_2023[11]), 
            .\SLO_buf[16]_adj_614 (SLO_buf_adj_8127[16]), .\SLO_buf[26]_adj_615 (SLO_buf_adj_8127[26]), 
            .\spi_data_out_r_39__N_4419[12] (spi_data_out_r_39__N_4419[12]), 
            .\spi_data_out_r_39__N_2023[10] (spi_data_out_r_39__N_2023[10]), 
            .\SLO_buf[15]_adj_616 (SLO_buf_adj_8127[15]), .\SLO_buf[25]_adj_617 (SLO_buf_adj_8127[25]), 
            .\spi_data_out_r_39__N_4419[11] (spi_data_out_r_39__N_4419[11]), 
            .\SLO_buf[24]_adj_618 (SLO_buf_adj_8127[24]), .\spi_data_out_r_39__N_4419[10] (spi_data_out_r_39__N_4419[10]), 
            .\SLO_buf[13]_adj_619 (SLO_buf_adj_8127[13]), .\SLO_buf[23]_adj_620 (SLO_buf_adj_8127[23]), 
            .\spi_data_out_r_39__N_4419[9] (spi_data_out_r_39__N_4419[9]), 
            .\SLO_buf[12]_adj_621 (SLO_buf_adj_8127[12]), .\SLO_buf[22]_adj_622 (SLO_buf_adj_8127[22]), 
            .\spi_data_out_r_39__N_4419[8] (spi_data_out_r_39__N_4419[8]), 
            .n25885(n25885), .n30087(n30087), .\quad_homing[1] (quad_homing_adj_7929[1]), 
            .n1(n1_adj_7669), .clk_enable_686(clk_enable_686), .clk_enable_260(clk_enable_260), 
            .clear_intrpt_adj_623(clear_intrpt), .intrpt_out_N_2642(intrpt_out_N_2642), 
            .intrpt_out_N_3068(intrpt_out_N_3068), .clk_enable_263(clk_enable_263), 
            .clk_enable_807(clk_enable_807), .n12467(n12467), .n20647(n20647), 
            .n18654(n18654), .n12435(n12435), .n26873(n26873), .clk_enable_320(clk_enable_320), 
            .n25877(n25877), .n30075(n30075), .\quad_homing[1]_adj_624 (quad_homing_adj_7777[1]), 
            .n1_adj_625(n1_adj_7668), .n30199(n30199), .n26821(n26821), 
            .clk_enable_684(clk_enable_684), .n26089(n26089), .n26091(n26091), 
            .clk_enable_255(clk_enable_255), .EM_STOP(EM_STOP), .clk_enable_23(clk_enable_23), 
            .n26947(n26947), .clk_enable_253(clk_enable_253), .pwm_out_N_3169(pwm_out_N_3169), 
            .pwm_out_N_3153(pwm_out_N_3153), .clk_enable_15(clk_enable_15), 
            .n26107(n26107), .n26113(n26113), .clear_intrpt_adj_626(clear_intrpt_adj_7665), 
            .intrpt_out_N_2997(intrpt_out_N_2997), .clk_enable_687(clk_enable_687), 
            .n30045(n30045), .clk_enable_759(clk_enable_759), .clk_enable_727(clk_enable_727), 
            .n11008(n11008), .pwm_out_1_N_6491(pwm_out_1_N_6491), .clk_enable_613(clk_enable_613), 
            .n26957(n26957), .clk_enable_520(clk_enable_520), .clk_enable_232(clk_enable_232), 
            .clk_enable_28(clk_enable_28), .clk_enable_226(clk_enable_226), 
            .clk_enable_639(clk_enable_639), .pwm_out_3_N_6530(pwm_out_3_N_6530), 
            .clk_enable_1105(clk_enable_1105), .pwm_out_4_N_6549(pwm_out_4_N_6549), 
            .clk_enable_1107(clk_enable_1107), .clk_enable_757(clk_enable_757), 
            .clk_enable_245(clk_enable_245), .pwm_out_2_N_6511(pwm_out_2_N_6511), 
            .clk_enable_22(clk_enable_22), .clk_enable_488(clk_enable_488), 
            .n26633(n26633), .clk_enable_641(clk_enable_641), .clk_enable_638(clk_enable_638), 
            .clk_enable_959(clk_enable_959), .clk_enable_235(clk_enable_235), 
            .intrpt_out_N_2713(intrpt_out_N_2713), .n57(n57), .reset_r_N_4129(reset_r_N_4129), 
            .clk_enable_761(clk_enable_761), .n29998(n29998), .clk_enable_738(clk_enable_738), 
            .n25881(n25881), .n30095(n30095), .\quad_homing[1]_adj_627 (quad_homing_adj_7815[1]), 
            .n1_adj_628(n1), .clk_enable_652(clk_enable_652), .quad_set_valid_N_2098(quad_set_valid_N_2098), 
            .clk_enable_683(clk_enable_683), .clk_enable_211(clk_enable_211), 
            .n2109(n2109), .n25893(n25893), .n30055(n30055), .\quad_homing[1]_adj_629 (quad_homing_adj_7891[1]), 
            .n1_adj_630(n1_adj_7712), .n25869(n25869), .n30043(n30043), 
            .\quad_homing[1]_adj_631 (quad_homing[1]), .n1_adj_632(n1_adj_7459), 
            .n25873(n25873), .n30091(n30091), .\quad_homing[1]_adj_633 (quad_homing_adj_7853[1]), 
            .n1_adj_634(n1_adj_7723), .n28476(n28476), .clk_enable_32(clk_enable_32), 
            .intrpt_out_N_2855(intrpt_out_N_2855), .clk_enable_178(clk_enable_178), 
            .intrpt_out_N_2784(intrpt_out_N_2784), .clk_enable_842(clk_enable_842), 
            .clk_enable_627(clk_enable_627), .clk_enable_234(clk_enable_234), 
            .quad_set_valid_N_2333(quad_set_valid_N_2333), .clk_enable_315(clk_enable_315), 
            .\SLO_buf[11]_adj_635 (SLO_buf_adj_8127[11]), .\SLO_buf[21]_adj_636 (SLO_buf_adj_8127[21]), 
            .\spi_data_out_r_39__N_4419[7] (spi_data_out_r_39__N_4419[7]), 
            .clk_enable_256(clk_enable_256), .n29999(n29999), .clk_enable_12(clk_enable_12), 
            .clk_enable_749(clk_enable_749), .clk_enable_388(clk_enable_388), 
            .n26207(n26207), .clk_enable_898(clk_enable_898), .clk_enable_180(clk_enable_180), 
            .n18_adj_637(n18), .n2193(n2193), .\SLO_buf[10]_adj_638 (SLO_buf_adj_8127[10]), 
            .\SLO_buf[20]_adj_639 (SLO_buf_adj_8127[20]), .\spi_data_out_r_39__N_4419[6] (spi_data_out_r_39__N_4419[6]), 
            .clk_enable_244(clk_enable_244), .intrpt_out_N_2926(intrpt_out_N_2926), 
            .pwm_out_1_N_6306(pwm_out_1_N_6306), .clk_100k_enable_1(clk_100k_enable_1), 
            .n25889(n25889), .n30083(n30083), .\quad_homing[1]_adj_640 (quad_homing_adj_7967[1]), 
            .n1_adj_641(n1_adj_7667), .clk_enable_595(clk_enable_595), .n30039(n30039), 
            .\spi_data_out_r_39__N_2023[9] (spi_data_out_r_39__N_2023[9]), 
            .\spi_data_out_r_39__N_1083[24] (spi_data_out_r_39__N_1083[24]), 
            .clear_intrpt_N_3001(clear_intrpt_N_3001), .\spi_data_out_r_39__N_2023[8] (spi_data_out_r_39__N_2023[8]), 
            .\spi_data_out_r_39__N_1083[11] (spi_data_out_r_39__N_1083[11]), 
            .\spi_data_out_r_39__N_2023[7] (spi_data_out_r_39__N_2023[7]), 
            .\spi_data_out_r_39__N_1083[27] (spi_data_out_r_39__N_1083[27]), 
            .\spi_data_out_r_39__N_4419[5] (spi_data_out_r_39__N_4419[5]), 
            .\spi_data_out_r_39__N_4419[4] (spi_data_out_r_39__N_4419[4]), 
            .\spi_data_out_r_39__N_2023[6] (spi_data_out_r_39__N_2023[6]), 
            .n27095(n27095), .spi_data_out_r_39__N_1868(spi_data_out_r_39__N_1868), 
            .n29992(n29992), .\spi_data_out_r_39__N_4419[3] (spi_data_out_r_39__N_4419[3]), 
            .\spi_data_out_r_39__N_2023[5] (spi_data_out_r_39__N_2023[5]), 
            .\spi_data_out_r_39__N_2023[24] (spi_data_out_r_39__N_2023[24]), 
            .\spi_data_out_r_39__N_4419[2] (spi_data_out_r_39__N_4419[2]), 
            .spi_data_out_r_39__N_5191(spi_data_out_r_39__N_5191), .spi_data_out_r_39__N_5534(spi_data_out_r_39__N_5534), 
            .spi_data_out_r_39__N_5877(spi_data_out_r_39__N_5877), .\spi_data_out_r_39__N_1083[23] (spi_data_out_r_39__N_1083[23]), 
            .spi_data_out_r_39__N_6220(spi_data_out_r_39__N_6220), .\spi_data_out_r_39__N_2023[4] (spi_data_out_r_39__N_2023[4]), 
            .\spi_data_out_r_39__N_2023[23] (spi_data_out_r_39__N_2023[23]), 
            .\spi_data_out_r_39__N_1083[1] (spi_data_out_r_39__N_1083[1]), 
            .\spi_data_out_r_39__N_1083[26] (spi_data_out_r_39__N_1083[26]), 
            .spi_data_out_r_39__N_1398(spi_data_out_r_39__N_1398), .\spi_data_out_r_39__N_1083[25] (spi_data_out_r_39__N_1083[25]), 
            .\spi_data_out_r_39__N_1083[30] (spi_data_out_r_39__N_1083[30]), 
            .n30013(n30013), .\spi_data_out_r_39__N_2023[3] (spi_data_out_r_39__N_2023[3]), 
            .\SLO_buf[5]_adj_642 (SLO_buf_adj_8127[5]), .\spi_data_out_r_39__N_4419[1] (spi_data_out_r_39__N_4419[1]), 
            .\spi_data_out_r_39__N_2023[2] (spi_data_out_r_39__N_2023[2]), 
            .\spi_data_out_r_39__N_2023[1] (spi_data_out_r_39__N_2023[1]), 
            .\spi_data_out_r_39__N_1083[10] (spi_data_out_r_39__N_1083[10]), 
            .\spi_data_out_r_39__N_2023[0] (spi_data_out_r_39__N_2023[0]), 
            .\spi_data_out_r_39__N_2023[22] (spi_data_out_r_39__N_2023[22]), 
            .n30007(n30007), .clk_enable_38(clk_enable_38), .\spi_data_out_r_39__N_2023[21] (spi_data_out_r_39__N_2023[21]), 
            .n30020(n30020), .\spi_data_out_r_39__N_2023[31] (spi_data_out_r_39__N_2023[31]), 
            .clk_enable_227(clk_enable_227), .\spi_data_out_r_39__N_2023[30] (spi_data_out_r_39__N_2023[30]), 
            .\spi_data_out_r_39__N_2023[29] (spi_data_out_r_39__N_2023[29]), 
            .\spi_data_out_r_39__N_1083[28] (spi_data_out_r_39__N_1083[28]), 
            .\spi_data_out_r_39__N_2023[28] (spi_data_out_r_39__N_2023[28]), 
            .\spi_data_out_r_39__N_2023[27] (spi_data_out_r_39__N_2023[27]), 
            .\spi_data_out_r_39__N_1083[21] (spi_data_out_r_39__N_1083[21]), 
            .n22554(n22554), .pwm(pwm), .n4_adj_643(n4), .\status_cntr[11] (status_cntr[11]), 
            .\spi_data_out_r_39__N_1083[0] (spi_data_out_r_39__N_1083[0]), 
            .spi_data_out_r_39__N_2103(spi_data_out_r_39__N_2103), .spi_data_out_r_39__N_1163(spi_data_out_r_39__N_1163), 
            .\spi_data_out_r_39__N_2493[0] (spi_data_out_r_39__N_2493[0]), 
            .\spi_data_out_r_39__N_2493[31] (spi_data_out_r_39__N_2493[31]), 
            .\spi_data_out_r_39__N_2493[30] (spi_data_out_r_39__N_2493[30]), 
            .spi_data_out_r_39__N_1633(spi_data_out_r_39__N_1633), .spi_data_out_r_39__N_2573(spi_data_out_r_39__N_2573)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(177[3] 197[2])
    \stepper(DEV_ID=1,UART_ADDRESS_WIDTH=4)  \stepper_ins_1..u_stepper  (.reset_r(reset_r_adj_7671), 
            .clk(clk), .clk_enable_12(clk_enable_12), .n30185(n30185), 
            .n29999(n29999), .clk_1MHz(clk_1MHz), .GND_net(GND_net), .resetn_c(resetn_c), 
            .pin_io_c_18(pin_io_c_18), .n30098(n30098), .spi_data_out_r_39__N_4168({spi_data_out_r_39__N_4168}), 
            .\spi_data_out_r_39__N_4419[0] (spi_data_out_r_39__N_4419[0]), 
            .clk_enable_759(clk_enable_759), .\spi_data_r[0] (spi_data_r[0]), 
            .\SLO_buf[0] (SLO_buf_adj_8127[0]), .n29992(n29992), .\SLO_buf[13] (SLO_buf_adj_8127[13]), 
            .\SLO_buf[12] (SLO_buf_adj_8127[12]), .\SLO_buf[11] (SLO_buf_adj_8127[11]), 
            .\SLO_buf[10] (SLO_buf_adj_8127[10]), .\spi_data_out_r_39__N_4419[35] (spi_data_out_r_39__N_4419[35]), 
            .\spi_data_out_r_39__N_4419[34] (spi_data_out_r_39__N_4419[34]), 
            .\spi_data_out_r_39__N_4419[33] (spi_data_out_r_39__N_4419[33]), 
            .\spi_data_out_r_39__N_4419[32] (spi_data_out_r_39__N_4419[32]), 
            .\spi_data_out_r_39__N_4419[15] (spi_data_out_r_39__N_4419[15]), 
            .\spi_data_out_r_39__N_4419[14] (spi_data_out_r_39__N_4419[14]), 
            .\spi_data_out_r_39__N_4419[13] (spi_data_out_r_39__N_4419[13]), 
            .\spi_data_out_r_39__N_4419[12] (spi_data_out_r_39__N_4419[12]), 
            .\spi_data_out_r_39__N_4419[11] (spi_data_out_r_39__N_4419[11]), 
            .\spi_data_out_r_39__N_4419[10] (spi_data_out_r_39__N_4419[10]), 
            .\spi_data_out_r_39__N_4419[9] (spi_data_out_r_39__N_4419[9]), 
            .\spi_data_out_r_39__N_4419[8] (spi_data_out_r_39__N_4419[8]), 
            .\spi_data_out_r_39__N_4419[7] (spi_data_out_r_39__N_4419[7]), 
            .\spi_data_out_r_39__N_4419[6] (spi_data_out_r_39__N_4419[6]), 
            .\spi_data_out_r_39__N_4419[5] (spi_data_out_r_39__N_4419[5]), 
            .\spi_data_out_r_39__N_4419[4] (spi_data_out_r_39__N_4419[4]), 
            .\spi_data_out_r_39__N_4419[3] (spi_data_out_r_39__N_4419[3]), 
            .\spi_data_out_r_39__N_4419[2] (spi_data_out_r_39__N_4419[2]), 
            .\spi_data_out_r_39__N_4419[1] (spi_data_out_r_39__N_4419[1]), 
            .\quad_homing[0] (quad_homing_adj_7777[0]), .pin_io_c_14(pin_io_c_14), 
            .n25877(n25877), .spi_data_out_r_39__N_4208(spi_data_out_r_39__N_4208), 
            .spi_data_out_r_39__N_4505(spi_data_out_r_39__N_4505), .digital_output_r(digital_output_r_adj_7672), 
            .clk_enable_256(clk_enable_256), .n28555(n28555), .\quad_a[1] (quad_a[1]), 
            .pin_io_out_19(pin_io_out_19), .\quad_b[1] (quad_b[1]), .uart_slot_en({uart_slot_en}), 
            .n30095(n30095), .n28(n28), .\spi_data_r[1] (spi_data_r[1]), 
            .\spi_data_r[2] (spi_data_r[2]), .\SLO_buf[1] (SLO_buf_adj_8127[1]), 
            .\SLO_buf[2] (SLO_buf_adj_8127[2]), .\SLO_buf[3] (SLO_buf_adj_8127[3]), 
            .\SLO_buf[4] (SLO_buf_adj_8127[4]), .\SLO_buf[5] (SLO_buf_adj_8127[5]), 
            .\SLO_buf[6] (SLO_buf_adj_8127[6]), .\SLO_buf[7] (SLO_buf_adj_8127[7]), 
            .\SLO_buf[8] (SLO_buf_adj_8127[8]), .\SLO_buf[9] (SLO_buf_adj_8127[9]), 
            .\SLO_buf[14] (SLO_buf_adj_8127[14]), .\SLO_buf[15] (SLO_buf_adj_8127[15]), 
            .\SLO_buf[16] (SLO_buf_adj_8127[16]), .\SLO_buf[17] (SLO_buf_adj_8127[17]), 
            .\SLO_buf[18] (SLO_buf_adj_8127[18]), .\SLO_buf[19] (SLO_buf_adj_8127[19]), 
            .\SLO_buf[20] (SLO_buf_adj_8127[20]), .\SLO_buf[21] (SLO_buf_adj_8127[21]), 
            .\SLO_buf[22] (SLO_buf_adj_8127[22]), .\SLO_buf[23] (SLO_buf_adj_8127[23]), 
            .\SLO_buf[24] (SLO_buf_adj_8127[24]), .\SLO_buf[25] (SLO_buf_adj_8127[25]), 
            .\SLO_buf[26] (SLO_buf_adj_8127[26]), .\SLO_buf[27] (SLO_buf_adj_8127[27]), 
            .\SLO_buf[28] (SLO_buf_adj_8127[28]), .\SLO_buf[29] (SLO_buf_adj_8127[29]), 
            .NSL(NSL_adj_7673), .UC_TXD0_c(UC_TXD0_c), .OW_ID_N_4461(OW_ID_N_4461), 
            .OW_ID_N_4467(OW_ID_N_4467), .n30050(n30050), .n30041(n30041), 
            .n30075(n30075), .pin_io_c_13(pin_io_c_13), .\pin_intrpt[4] (pin_intrpt[4]), 
            .pin_io_out_15(pin_io_out_15), .n29944(n29944), .pin_io_c_12(pin_io_c_12), 
            .\pin_intrpt[3] (pin_intrpt[3]), .\pin_intrpt[5] (pin_intrpt[5]), 
            .n7277(n7277), .ENC_O_N_4469(ENC_O_N_4469), .n30118(n30118), 
            .n30049(n30049), .\mode[2] (n31091[2]), .n9(n9_adj_7674)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(354[3] 397[2])
    \quad_decoder(DEV_ID=2)  \quad_ins_2..u_quad_decoder  (.quad_homing({quad_homing_adj_7815}), 
            .clk(clk), .clk_enable_488(clk_enable_488), .n30185(n30185), 
            .\spi_data_r[0] (spi_data_r[0]), .quad_count({quad_count_adj_7816}), 
            .\quad_b[2] (quad_b[2]), .\spi_data_out_r_39__N_1404[0] (spi_data_out_r_39__N_1404[0]), 
            .\spi_data_out_r_39__N_1553[0] (spi_data_out_r_39__N_1553[0]), 
            .quad_buffer({quad_buffer_adj_7817}), .\pin_intrpt[8] (pin_intrpt[8]), 
            .clk_enable_211(clk_enable_211), .\quad_a[2] (quad_a[2]), .\spi_data_r[31] (spi_data_r[31]), 
            .\spi_data_r[30] (spi_data_r[30]), .\spi_data_r[29] (spi_data_r[29]), 
            .\spi_data_r[28] (spi_data_r[28]), .\spi_data_r[27] (spi_data_r[27]), 
            .\spi_data_r[26] (spi_data_r[26]), .\spi_data_r[25] (spi_data_r[25]), 
            .\spi_data_r[24] (spi_data_r[24]), .\spi_data_r[23] (spi_data_r[23]), 
            .\spi_data_r[22] (spi_data_r[22]), .\spi_data_r[21] (spi_data_r[21]), 
            .\spi_data_r[20] (spi_data_r[20]), .\spi_data_r[19] (spi_data_r[19]), 
            .\spi_data_r[18] (spi_data_r[18]), .\spi_data_r[17] (spi_data_r[17]), 
            .\spi_data_r[16] (spi_data_r[16]), .\spi_data_r[15] (spi_data_r[15]), 
            .\spi_data_r[14] (spi_data_r[14]), .\spi_data_r[13] (spi_data_r[13]), 
            .\spi_data_r[12] (spi_data_r[12]), .\spi_data_r[11] (spi_data_r[11]), 
            .\spi_data_r[10] (spi_data_r[10]), .\spi_data_r[9] (spi_data_r[9]), 
            .\spi_data_r[8] (spi_data_r[8]), .\spi_data_r[7] (spi_data_r[7]), 
            .\spi_data_r[6] (spi_data_r[6]), .\spi_data_r[5] (spi_data_r[5]), 
            .\spi_data_r[4] (spi_data_r[4]), .\spi_data_r[3] (spi_data_r[3]), 
            .\spi_data_r[2] (spi_data_r[2]), .\spi_data_r[1] (spi_data_r[1]), 
            .spi_data_out_r_39__N_1444(spi_data_out_r_39__N_1444), .spi_data_out_r_39__N_1633(spi_data_out_r_39__N_1633), 
            .n29993(n29993), .\spi_data_out_r_39__N_1404[31] (spi_data_out_r_39__N_1404[31]), 
            .\spi_data_out_r_39__N_1553[31] (spi_data_out_r_39__N_1553[31]), 
            .\spi_data_out_r_39__N_1404[30] (spi_data_out_r_39__N_1404[30]), 
            .\spi_data_out_r_39__N_1553[30] (spi_data_out_r_39__N_1553[30]), 
            .\spi_data_out_r_39__N_1404[29] (spi_data_out_r_39__N_1404[29]), 
            .\spi_data_out_r_39__N_1553[29] (spi_data_out_r_39__N_1553[29]), 
            .\spi_data_out_r_39__N_1404[28] (spi_data_out_r_39__N_1404[28]), 
            .\spi_data_out_r_39__N_1553[28] (spi_data_out_r_39__N_1553[28]), 
            .\spi_data_out_r_39__N_1404[27] (spi_data_out_r_39__N_1404[27]), 
            .\spi_data_out_r_39__N_1553[27] (spi_data_out_r_39__N_1553[27]), 
            .\spi_data_out_r_39__N_1404[26] (spi_data_out_r_39__N_1404[26]), 
            .\spi_data_out_r_39__N_1553[26] (spi_data_out_r_39__N_1553[26]), 
            .\spi_data_out_r_39__N_1404[25] (spi_data_out_r_39__N_1404[25]), 
            .\spi_data_out_r_39__N_1553[25] (spi_data_out_r_39__N_1553[25]), 
            .\spi_data_out_r_39__N_1404[24] (spi_data_out_r_39__N_1404[24]), 
            .\spi_data_out_r_39__N_1553[24] (spi_data_out_r_39__N_1553[24]), 
            .\spi_data_out_r_39__N_1404[23] (spi_data_out_r_39__N_1404[23]), 
            .\spi_data_out_r_39__N_1553[23] (spi_data_out_r_39__N_1553[23]), 
            .\spi_data_out_r_39__N_1404[22] (spi_data_out_r_39__N_1404[22]), 
            .\spi_data_out_r_39__N_1553[22] (spi_data_out_r_39__N_1553[22]), 
            .\spi_data_out_r_39__N_1404[21] (spi_data_out_r_39__N_1404[21]), 
            .\spi_data_out_r_39__N_1553[21] (spi_data_out_r_39__N_1553[21]), 
            .\spi_data_out_r_39__N_1404[20] (spi_data_out_r_39__N_1404[20]), 
            .\spi_data_out_r_39__N_1553[20] (spi_data_out_r_39__N_1553[20]), 
            .\spi_data_out_r_39__N_1404[19] (spi_data_out_r_39__N_1404[19]), 
            .\spi_data_out_r_39__N_1553[19] (spi_data_out_r_39__N_1553[19]), 
            .\spi_data_out_r_39__N_1404[18] (spi_data_out_r_39__N_1404[18]), 
            .\spi_data_out_r_39__N_1553[18] (spi_data_out_r_39__N_1553[18]), 
            .\spi_data_out_r_39__N_1404[17] (spi_data_out_r_39__N_1404[17]), 
            .\spi_data_out_r_39__N_1553[17] (spi_data_out_r_39__N_1553[17]), 
            .\spi_data_out_r_39__N_1404[16] (spi_data_out_r_39__N_1404[16]), 
            .\spi_data_out_r_39__N_1553[16] (spi_data_out_r_39__N_1553[16]), 
            .\spi_data_out_r_39__N_1404[15] (spi_data_out_r_39__N_1404[15]), 
            .\spi_data_out_r_39__N_1553[15] (spi_data_out_r_39__N_1553[15]), 
            .\spi_data_out_r_39__N_1404[14] (spi_data_out_r_39__N_1404[14]), 
            .\spi_data_out_r_39__N_1553[14] (spi_data_out_r_39__N_1553[14]), 
            .\spi_data_out_r_39__N_1404[13] (spi_data_out_r_39__N_1404[13]), 
            .\spi_data_out_r_39__N_1553[13] (spi_data_out_r_39__N_1553[13]), 
            .\spi_data_out_r_39__N_1404[12] (spi_data_out_r_39__N_1404[12]), 
            .\spi_data_out_r_39__N_1553[12] (spi_data_out_r_39__N_1553[12]), 
            .\spi_data_out_r_39__N_1404[11] (spi_data_out_r_39__N_1404[11]), 
            .\spi_data_out_r_39__N_1553[11] (spi_data_out_r_39__N_1553[11]), 
            .\spi_data_out_r_39__N_1404[10] (spi_data_out_r_39__N_1404[10]), 
            .\spi_data_out_r_39__N_1553[10] (spi_data_out_r_39__N_1553[10]), 
            .\spi_data_out_r_39__N_1404[9] (spi_data_out_r_39__N_1404[9]), 
            .\spi_data_out_r_39__N_1553[9] (spi_data_out_r_39__N_1553[9]), 
            .\spi_data_out_r_39__N_1404[8] (spi_data_out_r_39__N_1404[8]), 
            .\spi_data_out_r_39__N_1553[8] (spi_data_out_r_39__N_1553[8]), 
            .\spi_data_out_r_39__N_1404[7] (spi_data_out_r_39__N_1404[7]), 
            .\spi_data_out_r_39__N_1553[7] (spi_data_out_r_39__N_1553[7]), 
            .\spi_data_out_r_39__N_1404[6] (spi_data_out_r_39__N_1404[6]), 
            .\spi_data_out_r_39__N_1553[6] (spi_data_out_r_39__N_1553[6]), 
            .\spi_data_out_r_39__N_1404[5] (spi_data_out_r_39__N_1404[5]), 
            .\spi_data_out_r_39__N_1553[5] (spi_data_out_r_39__N_1553[5]), 
            .\spi_data_out_r_39__N_1404[4] (spi_data_out_r_39__N_1404[4]), 
            .\spi_data_out_r_39__N_1553[4] (spi_data_out_r_39__N_1553[4]), 
            .\spi_data_out_r_39__N_1404[3] (spi_data_out_r_39__N_1404[3]), 
            .\spi_data_out_r_39__N_1553[3] (spi_data_out_r_39__N_1553[3]), 
            .\spi_data_out_r_39__N_1404[2] (spi_data_out_r_39__N_1404[2]), 
            .\spi_data_out_r_39__N_1553[2] (spi_data_out_r_39__N_1553[2]), 
            .\spi_data_out_r_39__N_1404[1] (spi_data_out_r_39__N_1404[1]), 
            .\spi_data_out_r_39__N_1553[1] (spi_data_out_r_39__N_1553[1]), 
            .resetn_c(resetn_c), .n1(n1), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(263[3] 283[2])
    quad_decoder \quad_ins_0..u_quad_decoder  (.quad_count({quad_count}), 
            .clk(clk), .n30185(n30185), .\quad_b[0] (quad_b[0]), .\spi_data_out_r_39__N_934[0] (spi_data_out_r_39__N_934[0]), 
            .\spi_data_out_r_39__N_1083[0] (spi_data_out_r_39__N_1083[0]), 
            .quad_buffer({quad_buffer}), .\pin_intrpt[2] (pin_intrpt[2]), 
            .quad_set_valid_N_1158(quad_set_valid_N_1158), .\quad_a[0] (quad_a[0]), 
            .quad_homing({quad_homing}), .clk_enable_757(clk_enable_757), 
            .\spi_data_r[0] (spi_data_r[0]), .clk_enable_807(clk_enable_807), 
            .GND_net(GND_net), .spi_data_out_r_39__N_974(spi_data_out_r_39__N_974), 
            .spi_data_out_r_39__N_1163(spi_data_out_r_39__N_1163), .\spi_cmd_r[2] (spi_cmd_r[2]), 
            .\spi_addr_r[7] (spi_addr_r[7]), .n28328(n28328), .\spi_data_out_r_39__N_934[31] (spi_data_out_r_39__N_934[31]), 
            .\spi_data_out_r_39__N_1083[31] (spi_data_out_r_39__N_1083[31]), 
            .\spi_data_out_r_39__N_934[30] (spi_data_out_r_39__N_934[30]), 
            .\spi_data_out_r_39__N_1083[30] (spi_data_out_r_39__N_1083[30]), 
            .\spi_data_out_r_39__N_934[29] (spi_data_out_r_39__N_934[29]), 
            .\spi_data_out_r_39__N_1083[29] (spi_data_out_r_39__N_1083[29]), 
            .\spi_data_out_r_39__N_934[28] (spi_data_out_r_39__N_934[28]), 
            .\spi_data_out_r_39__N_1083[28] (spi_data_out_r_39__N_1083[28]), 
            .\spi_data_out_r_39__N_934[27] (spi_data_out_r_39__N_934[27]), 
            .\spi_data_out_r_39__N_1083[27] (spi_data_out_r_39__N_1083[27]), 
            .\spi_data_out_r_39__N_934[26] (spi_data_out_r_39__N_934[26]), 
            .\spi_data_out_r_39__N_1083[26] (spi_data_out_r_39__N_1083[26]), 
            .\spi_data_out_r_39__N_934[25] (spi_data_out_r_39__N_934[25]), 
            .\spi_data_out_r_39__N_1083[25] (spi_data_out_r_39__N_1083[25]), 
            .\spi_data_out_r_39__N_934[24] (spi_data_out_r_39__N_934[24]), 
            .\spi_data_out_r_39__N_1083[24] (spi_data_out_r_39__N_1083[24]), 
            .\spi_data_out_r_39__N_934[23] (spi_data_out_r_39__N_934[23]), 
            .\spi_data_out_r_39__N_1083[23] (spi_data_out_r_39__N_1083[23]), 
            .\spi_data_out_r_39__N_934[22] (spi_data_out_r_39__N_934[22]), 
            .\spi_data_out_r_39__N_1083[22] (spi_data_out_r_39__N_1083[22]), 
            .\spi_data_out_r_39__N_934[21] (spi_data_out_r_39__N_934[21]), 
            .\spi_data_out_r_39__N_1083[21] (spi_data_out_r_39__N_1083[21]), 
            .\spi_data_out_r_39__N_934[20] (spi_data_out_r_39__N_934[20]), 
            .\spi_data_out_r_39__N_1083[20] (spi_data_out_r_39__N_1083[20]), 
            .\spi_data_out_r_39__N_934[19] (spi_data_out_r_39__N_934[19]), 
            .\spi_data_out_r_39__N_1083[19] (spi_data_out_r_39__N_1083[19]), 
            .\spi_data_out_r_39__N_934[18] (spi_data_out_r_39__N_934[18]), 
            .\spi_data_out_r_39__N_1083[18] (spi_data_out_r_39__N_1083[18]), 
            .\spi_data_out_r_39__N_934[17] (spi_data_out_r_39__N_934[17]), 
            .\spi_data_out_r_39__N_1083[17] (spi_data_out_r_39__N_1083[17]), 
            .\spi_data_out_r_39__N_934[16] (spi_data_out_r_39__N_934[16]), 
            .\spi_data_out_r_39__N_1083[16] (spi_data_out_r_39__N_1083[16]), 
            .\spi_data_out_r_39__N_934[15] (spi_data_out_r_39__N_934[15]), 
            .\spi_data_out_r_39__N_1083[15] (spi_data_out_r_39__N_1083[15]), 
            .\spi_data_out_r_39__N_934[14] (spi_data_out_r_39__N_934[14]), 
            .\spi_data_out_r_39__N_1083[14] (spi_data_out_r_39__N_1083[14]), 
            .\spi_data_out_r_39__N_934[13] (spi_data_out_r_39__N_934[13]), 
            .\spi_data_out_r_39__N_1083[13] (spi_data_out_r_39__N_1083[13]), 
            .\spi_data_out_r_39__N_934[12] (spi_data_out_r_39__N_934[12]), 
            .\spi_data_out_r_39__N_1083[12] (spi_data_out_r_39__N_1083[12]), 
            .\spi_data_out_r_39__N_934[11] (spi_data_out_r_39__N_934[11]), 
            .\spi_data_out_r_39__N_1083[11] (spi_data_out_r_39__N_1083[11]), 
            .\spi_data_out_r_39__N_934[10] (spi_data_out_r_39__N_934[10]), 
            .\spi_data_out_r_39__N_1083[10] (spi_data_out_r_39__N_1083[10]), 
            .\spi_data_out_r_39__N_934[9] (spi_data_out_r_39__N_934[9]), .\spi_data_out_r_39__N_1083[9] (spi_data_out_r_39__N_1083[9]), 
            .\spi_data_out_r_39__N_934[8] (spi_data_out_r_39__N_934[8]), .\spi_data_out_r_39__N_1083[8] (spi_data_out_r_39__N_1083[8]), 
            .\spi_data_out_r_39__N_934[7] (spi_data_out_r_39__N_934[7]), .\spi_data_out_r_39__N_1083[7] (spi_data_out_r_39__N_1083[7]), 
            .\spi_data_out_r_39__N_934[6] (spi_data_out_r_39__N_934[6]), .\spi_data_out_r_39__N_1083[6] (spi_data_out_r_39__N_1083[6]), 
            .\spi_data_out_r_39__N_934[5] (spi_data_out_r_39__N_934[5]), .\spi_data_out_r_39__N_1083[5] (spi_data_out_r_39__N_1083[5]), 
            .\spi_data_out_r_39__N_934[4] (spi_data_out_r_39__N_934[4]), .\spi_data_out_r_39__N_1083[4] (spi_data_out_r_39__N_1083[4]), 
            .\spi_data_out_r_39__N_934[3] (spi_data_out_r_39__N_934[3]), .\spi_data_out_r_39__N_1083[3] (spi_data_out_r_39__N_1083[3]), 
            .\spi_data_out_r_39__N_934[2] (spi_data_out_r_39__N_934[2]), .\spi_data_out_r_39__N_1083[2] (spi_data_out_r_39__N_1083[2]), 
            .\spi_data_out_r_39__N_934[1] (spi_data_out_r_39__N_934[1]), .\spi_data_out_r_39__N_1083[1] (spi_data_out_r_39__N_1083[1]), 
            .\spi_data_r[1] (spi_data_r[1]), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[3] (spi_data_r[3]), .\spi_data_r[4] (spi_data_r[4]), 
            .\spi_data_r[5] (spi_data_r[5]), .\spi_data_r[6] (spi_data_r[6]), 
            .\spi_data_r[7] (spi_data_r[7]), .\spi_data_r[8] (spi_data_r[8]), 
            .\spi_data_r[9] (spi_data_r[9]), .\spi_data_r[10] (spi_data_r[10]), 
            .\spi_data_r[11] (spi_data_r[11]), .\spi_data_r[12] (spi_data_r[12]), 
            .\spi_data_r[13] (spi_data_r[13]), .\spi_data_r[14] (spi_data_r[14]), 
            .\spi_data_r[15] (spi_data_r[15]), .\spi_data_r[16] (spi_data_r[16]), 
            .\spi_data_r[17] (spi_data_r[17]), .\spi_data_r[18] (spi_data_r[18]), 
            .\spi_data_r[19] (spi_data_r[19]), .\spi_data_r[20] (spi_data_r[20]), 
            .\spi_data_r[21] (spi_data_r[21]), .\spi_data_r[22] (spi_data_r[22]), 
            .\spi_data_r[23] (spi_data_r[23]), .\spi_data_r[24] (spi_data_r[24]), 
            .\spi_data_r[25] (spi_data_r[25]), .\spi_data_r[26] (spi_data_r[26]), 
            .\spi_data_r[27] (spi_data_r[27]), .\spi_data_r[28] (spi_data_r[28]), 
            .\spi_data_r[29] (spi_data_r[29]), .\spi_data_r[30] (spi_data_r[30]), 
            .\spi_data_r[31] (spi_data_r[31]), .n28340(n28340), .n23916(n23916), 
            .n26327(n26327), .quad_set_valid_N_2098(quad_set_valid_N_2098), 
            .\spi_addr_r[6] (spi_addr_r[6]), .n30209(n30209), .n28384(n28384), 
            .\spi_addr_r[2] (spi_addr_r[2]), .n28524(n28524), .n24169(n24169), 
            .\spi_addr_r[0] (spi_addr_r[0]), .\spi_addr_r[1] (spi_addr_r[1]), 
            .reset_r_N_4129(reset_r_N_4129), .n1(n1_adj_7459), .resetn_c(resetn_c), 
            .n25547(n25547)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(263[3] 283[2])
    \stepper(DEV_ID=6,UART_ADDRESS_WIDTH=4)  \stepper_ins_6..u_stepper  (.\spi_data_out_r_39__N_5540[4] (spi_data_out_r_39__N_5540[4]), 
            .spi_data_out_r_39__N_5580(spi_data_out_r_39__N_5580), .\spi_data_out_r_39__N_4511[4] (spi_data_out_r_39__N_4511[4]), 
            .spi_data_out_r_39__N_4551(spi_data_out_r_39__N_4551), .clk(clk), 
            .\spi_data_out_r_39__N_1404[4] (spi_data_out_r_39__N_1404[4]), 
            .\spi_data_out_r_39__N_1639[4] (spi_data_out_r_39__N_1639[4]), 
            .spi_data_out_r_39__N_1444(spi_data_out_r_39__N_1444), .spi_data_out_r_39__N_1679(spi_data_out_r_39__N_1679), 
            .\spi_data_out_r_39__N_1874[4] (spi_data_out_r_39__N_1874[4]), 
            .spi_data_out_r_39__N_1914(spi_data_out_r_39__N_1914), .\spi_data_out_r_39__N_1169[4] (spi_data_out_r_39__N_1169[4]), 
            .spi_data_out_r_39__N_1209(spi_data_out_r_39__N_1209), .\spi_data_out_r_39__N_2109[4] (spi_data_out_r_39__N_2109[4]), 
            .\spi_data_out_r_39__N_934[4] (spi_data_out_r_39__N_934[4]), .spi_data_out_r_39__N_2149(spi_data_out_r_39__N_2149), 
            .spi_data_out_r_39__N_974(spi_data_out_r_39__N_974), .\spi_data_out_r_39__N_2344[4] (spi_data_out_r_39__N_2344[4]), 
            .spi_data_out_r_39__N_2384(spi_data_out_r_39__N_2384), .\spi_data_out_r_39__N_5197[4] (spi_data_out_r_39__N_5197[4]), 
            .\spi_data_out_r_39__N_4854[4] (spi_data_out_r_39__N_4854[4]), 
            .spi_data_out_r_39__N_5237(spi_data_out_r_39__N_5237), .spi_data_out_r_39__N_4894(spi_data_out_r_39__N_4894), 
            .spi_data_out_r_39__N_5923(spi_data_out_r_39__N_5923), .\spi_data_out_r[5] (spi_data_out_r[5]), 
            .\spi_data_out_r_39__N_3825[5] (spi_data_out_r_39__N_3825[5]), 
            .\spi_data_out_r_39__N_4168[5] (spi_data_out_r_39__N_4168[5]), 
            .spi_data_out_r_39__N_3865(spi_data_out_r_39__N_3865), .spi_data_out_r_39__N_4208(spi_data_out_r_39__N_4208), 
            .\spi_data_out_r_39__N_5540[5] (spi_data_out_r_39__N_5540[5]), 
            .reset_r(reset_r_adj_7720), .n30185(n30185), .n30028(n30028), 
            .NSL(NSL_adj_7722), .clk_1MHz(clk_1MHz), .\spi_data_out_r_39__N_4511[5] (spi_data_out_r_39__N_4511[5]), 
            .\spi_data_out_r_39__N_1404[5] (spi_data_out_r_39__N_1404[5]), 
            .\spi_data_out_r_39__N_1639[5] (spi_data_out_r_39__N_1639[5]), 
            .\spi_data_out_r_39__N_1874[5] (spi_data_out_r_39__N_1874[5]), 
            .\spi_data_out_r_39__N_1169[5] (spi_data_out_r_39__N_1169[5]), 
            .\spi_data_out_r_39__N_2109[5] (spi_data_out_r_39__N_2109[5]), 
            .\spi_data_out_r_39__N_934[5] (spi_data_out_r_39__N_934[5]), .\spi_data_out_r_39__N_2344[5] (spi_data_out_r_39__N_2344[5]), 
            .\spi_data_out_r_39__N_5197[5] (spi_data_out_r_39__N_5197[5]), 
            .\spi_data_out_r_39__N_4854[5] (spi_data_out_r_39__N_4854[5]), 
            .clk_enable_180(clk_enable_180), .\spi_data_r[0] (spi_data_r[0]), 
            .\spi_data_out_r[6] (spi_data_out_r[6]), .\spi_data_out_r_39__N_3825[6] (spi_data_out_r_39__N_3825[6]), 
            .\spi_data_out_r_39__N_4168[6] (spi_data_out_r_39__N_4168[6]), 
            .\spi_data_out_r_39__N_5540[6] (spi_data_out_r_39__N_5540[6]), 
            .\spi_data_out_r_39__N_4511[6] (spi_data_out_r_39__N_4511[6]), 
            .\spi_data_out_r_39__N_1404[6] (spi_data_out_r_39__N_1404[6]), 
            .\spi_data_out_r_39__N_1639[6] (spi_data_out_r_39__N_1639[6]), 
            .\spi_data_out_r_39__N_1874[6] (spi_data_out_r_39__N_1874[6]), 
            .\spi_data_out_r_39__N_1169[6] (spi_data_out_r_39__N_1169[6]), 
            .\spi_data_out_r_39__N_2109[6] (spi_data_out_r_39__N_2109[6]), 
            .\spi_data_out_r_39__N_934[6] (spi_data_out_r_39__N_934[6]), .\spi_data_out_r_39__N_2344[6] (spi_data_out_r_39__N_2344[6]), 
            .\spi_data_out_r_39__N_5197[6] (spi_data_out_r_39__N_5197[6]), 
            .\spi_data_out_r_39__N_4854[6] (spi_data_out_r_39__N_4854[6]), 
            .\spi_data_out_r[7] (spi_data_out_r[7]), .\spi_data_out_r_39__N_3825[7] (spi_data_out_r_39__N_3825[7]), 
            .\spi_data_out_r_39__N_4168[7] (spi_data_out_r_39__N_4168[7]), 
            .\spi_data_out_r_39__N_5540[7] (spi_data_out_r_39__N_5540[7]), 
            .\spi_data_out_r_39__N_4511[7] (spi_data_out_r_39__N_4511[7]), 
            .\spi_data_out_r_39__N_1404[7] (spi_data_out_r_39__N_1404[7]), 
            .\spi_data_out_r_39__N_1639[7] (spi_data_out_r_39__N_1639[7]), 
            .n30143(n30143), .\spi_data_out_r_39__N_1874[7] (spi_data_out_r_39__N_1874[7]), 
            .\spi_data_out_r_39__N_1169[7] (spi_data_out_r_39__N_1169[7]), 
            .\spi_data_out_r_39__N_2109[7] (spi_data_out_r_39__N_2109[7]), 
            .\spi_data_out_r_39__N_934[7] (spi_data_out_r_39__N_934[7]), .\spi_data_out_r_39__N_2344[7] (spi_data_out_r_39__N_2344[7]), 
            .\spi_data_out_r_39__N_5197[7] (spi_data_out_r_39__N_5197[7]), 
            .\spi_data_out_r_39__N_4854[7] (spi_data_out_r_39__N_4854[7]), 
            .resetn_c(resetn_c), .\spi_data_out_r[10] (spi_data_out_r[10]), 
            .\spi_data_out_r_39__N_3825[10] (spi_data_out_r_39__N_3825[10]), 
            .\spi_data_out_r_39__N_4168[10] (spi_data_out_r_39__N_4168[10]), 
            .\spi_data_r[2] (spi_data_r[2]), .\spi_data_r[1] (spi_data_r[1]), 
            .\spi_data_out_r_39__N_5540[10] (spi_data_out_r_39__N_5540[10]), 
            .\spi_data_out_r_39__N_4511[10] (spi_data_out_r_39__N_4511[10]), 
            .\spi_data_out_r_39__N_1404[10] (spi_data_out_r_39__N_1404[10]), 
            .\spi_data_out_r_39__N_1639[10] (spi_data_out_r_39__N_1639[10]), 
            .\spi_data_out_r_39__N_1874[10] (spi_data_out_r_39__N_1874[10]), 
            .\spi_data_out_r_39__N_1169[10] (spi_data_out_r_39__N_1169[10]), 
            .\spi_data_out_r_39__N_2109[10] (spi_data_out_r_39__N_2109[10]), 
            .\spi_data_out_r_39__N_934[10] (spi_data_out_r_39__N_934[10]), 
            .\spi_data_out_r_39__N_2344[10] (spi_data_out_r_39__N_2344[10]), 
            .\spi_data_out_r_39__N_5197[10] (spi_data_out_r_39__N_5197[10]), 
            .\spi_data_out_r_39__N_4854[10] (spi_data_out_r_39__N_4854[10]), 
            .\spi_data_out_r[11] (spi_data_out_r[11]), .\spi_data_out_r_39__N_3825[11] (spi_data_out_r_39__N_3825[11]), 
            .\spi_data_out_r_39__N_4168[11] (spi_data_out_r_39__N_4168[11]), 
            .\spi_data_out_r_39__N_5540[11] (spi_data_out_r_39__N_5540[11]), 
            .\spi_data_out_r_39__N_4511[11] (spi_data_out_r_39__N_4511[11]), 
            .\spi_data_out_r_39__N_1404[11] (spi_data_out_r_39__N_1404[11]), 
            .\spi_data_out_r_39__N_1639[11] (spi_data_out_r_39__N_1639[11]), 
            .\spi_data_out_r_39__N_1874[11] (spi_data_out_r_39__N_1874[11]), 
            .\spi_data_out_r_39__N_1169[11] (spi_data_out_r_39__N_1169[11]), 
            .\spi_data_out_r_39__N_2109[11] (spi_data_out_r_39__N_2109[11]), 
            .\spi_data_out_r_39__N_934[11] (spi_data_out_r_39__N_934[11]), 
            .\spi_data_out_r_39__N_2344[11] (spi_data_out_r_39__N_2344[11]), 
            .\spi_data_out_r_39__N_5197[11] (spi_data_out_r_39__N_5197[11]), 
            .\spi_data_out_r_39__N_4854[11] (spi_data_out_r_39__N_4854[11]), 
            .\spi_data_out_r[12] (spi_data_out_r[12]), .\spi_data_out_r_39__N_3825[12] (spi_data_out_r_39__N_3825[12]), 
            .\spi_data_out_r_39__N_4168[12] (spi_data_out_r_39__N_4168[12]), 
            .\spi_data_out_r_39__N_5540[12] (spi_data_out_r_39__N_5540[12]), 
            .\spi_data_out_r_39__N_4511[12] (spi_data_out_r_39__N_4511[12]), 
            .\spi_data_out_r_39__N_1404[12] (spi_data_out_r_39__N_1404[12]), 
            .\spi_data_out_r_39__N_1639[12] (spi_data_out_r_39__N_1639[12]), 
            .\spi_data_out_r_39__N_1874[12] (spi_data_out_r_39__N_1874[12]), 
            .\spi_data_out_r_39__N_1169[12] (spi_data_out_r_39__N_1169[12]), 
            .\spi_data_out_r_39__N_2109[12] (spi_data_out_r_39__N_2109[12]), 
            .\spi_data_out_r_39__N_934[12] (spi_data_out_r_39__N_934[12]), 
            .\spi_data_out_r_39__N_2344[12] (spi_data_out_r_39__N_2344[12]), 
            .\spi_data_out_r_39__N_5197[12] (spi_data_out_r_39__N_5197[12]), 
            .\spi_data_out_r_39__N_4854[12] (spi_data_out_r_39__N_4854[12]), 
            .\spi_data_out_r[13] (spi_data_out_r[13]), .\spi_data_out_r_39__N_3825[13] (spi_data_out_r_39__N_3825[13]), 
            .\spi_data_out_r_39__N_4168[13] (spi_data_out_r_39__N_4168[13]), 
            .digital_output_r(digital_output_r_adj_7721), .clk_enable_222(clk_enable_222), 
            .n28550(n28550), .\spi_data_out_r_39__N_5540[13] (spi_data_out_r_39__N_5540[13]), 
            .EM_STOP(EM_STOP), .n25741(n25741), .n23916(n23916), .\spi_data_out_r_39__N_4511[13] (spi_data_out_r_39__N_4511[13]), 
            .\spi_data_out_r_39__N_1404[13] (spi_data_out_r_39__N_1404[13]), 
            .\spi_data_out_r_39__N_1639[13] (spi_data_out_r_39__N_1639[13]), 
            .\spi_data_out_r_39__N_1874[13] (spi_data_out_r_39__N_1874[13]), 
            .\spi_data_out_r_39__N_1169[13] (spi_data_out_r_39__N_1169[13]), 
            .\spi_data_out_r_39__N_2109[13] (spi_data_out_r_39__N_2109[13]), 
            .\spi_data_out_r_39__N_934[13] (spi_data_out_r_39__N_934[13]), 
            .\spi_data_out_r_39__N_2344[13] (spi_data_out_r_39__N_2344[13]), 
            .\spi_data_out_r_39__N_5197[13] (spi_data_out_r_39__N_5197[13]), 
            .\spi_data_out_r_39__N_4854[13] (spi_data_out_r_39__N_4854[13]), 
            .\spi_data_out_r[14] (spi_data_out_r[14]), .\spi_data_out_r_39__N_3825[14] (spi_data_out_r_39__N_3825[14]), 
            .\spi_data_out_r_39__N_4168[14] (spi_data_out_r_39__N_4168[14]), 
            .\spi_data_out_r_39__N_5540[14] (spi_data_out_r_39__N_5540[14]), 
            .\spi_data_out_r_39__N_4511[14] (spi_data_out_r_39__N_4511[14]), 
            .\spi_data_out_r_39__N_1404[14] (spi_data_out_r_39__N_1404[14]), 
            .\spi_data_out_r_39__N_1639[14] (spi_data_out_r_39__N_1639[14]), 
            .\spi_data_out_r_39__N_1874[14] (spi_data_out_r_39__N_1874[14]), 
            .\spi_data_out_r_39__N_1169[14] (spi_data_out_r_39__N_1169[14]), 
            .\spi_data_out_r_39__N_2109[14] (spi_data_out_r_39__N_2109[14]), 
            .\spi_data_out_r_39__N_934[14] (spi_data_out_r_39__N_934[14]), 
            .\spi_data_out_r_39__N_2344[14] (spi_data_out_r_39__N_2344[14]), 
            .\spi_data_out_r_39__N_5197[14] (spi_data_out_r_39__N_5197[14]), 
            .\spi_data_out_r_39__N_4854[14] (spi_data_out_r_39__N_4854[14]), 
            .\spi_data_out_r[15] (spi_data_out_r[15]), .\spi_data_out_r_39__N_3825[15] (spi_data_out_r_39__N_3825[15]), 
            .\spi_data_out_r_39__N_4168[15] (spi_data_out_r_39__N_4168[15]), 
            .\spi_data_out_r_39__N_5540[15] (spi_data_out_r_39__N_5540[15]), 
            .\spi_data_out_r_39__N_4511[15] (spi_data_out_r_39__N_4511[15]), 
            .\spi_data_out_r_39__N_1404[15] (spi_data_out_r_39__N_1404[15]), 
            .\spi_data_out_r_39__N_1639[15] (spi_data_out_r_39__N_1639[15]), 
            .\spi_data_out_r_39__N_1874[15] (spi_data_out_r_39__N_1874[15]), 
            .\spi_data_out_r_39__N_1169[15] (spi_data_out_r_39__N_1169[15]), 
            .\spi_data_out_r_39__N_2109[15] (spi_data_out_r_39__N_2109[15]), 
            .\spi_data_out_r_39__N_934[15] (spi_data_out_r_39__N_934[15]), 
            .\spi_data_out_r_39__N_2344[15] (spi_data_out_r_39__N_2344[15]), 
            .\spi_data_out_r_39__N_5197[15] (spi_data_out_r_39__N_5197[15]), 
            .\spi_data_out_r_39__N_4854[15] (spi_data_out_r_39__N_4854[15]), 
            .\spi_data_out_r[16] (spi_data_out_r[16]), .\spi_data_out_r_39__N_3825[16] (spi_data_out_r_39__N_3825[16]), 
            .\spi_data_out_r_39__N_4168[16] (spi_data_out_r_39__N_4168[16]), 
            .\spi_data_out_r_39__N_5540[16] (spi_data_out_r_39__N_5540[16]), 
            .\spi_data_out_r_39__N_4511[16] (spi_data_out_r_39__N_4511[16]), 
            .\spi_data_out_r_39__N_1404[16] (spi_data_out_r_39__N_1404[16]), 
            .\spi_data_out_r_39__N_1639[16] (spi_data_out_r_39__N_1639[16]), 
            .\spi_data_out_r_39__N_1874[16] (spi_data_out_r_39__N_1874[16]), 
            .\spi_data_out_r_39__N_1169[16] (spi_data_out_r_39__N_1169[16]), 
            .\spi_data_out_r_39__N_2109[16] (spi_data_out_r_39__N_2109[16]), 
            .\spi_data_out_r_39__N_934[16] (spi_data_out_r_39__N_934[16]), 
            .\spi_data_out_r_39__N_2344[16] (spi_data_out_r_39__N_2344[16]), 
            .\spi_data_out_r_39__N_5197[16] (spi_data_out_r_39__N_5197[16]), 
            .\spi_data_out_r_39__N_4854[16] (spi_data_out_r_39__N_4854[16]), 
            .\spi_data_out_r[17] (spi_data_out_r[17]), .\spi_data_out_r_39__N_3825[17] (spi_data_out_r_39__N_3825[17]), 
            .\spi_data_out_r_39__N_4168[17] (spi_data_out_r_39__N_4168[17]), 
            .\spi_data_out_r_39__N_5540[17] (spi_data_out_r_39__N_5540[17]), 
            .\spi_data_out_r_39__N_4511[17] (spi_data_out_r_39__N_4511[17]), 
            .\spi_data_out_r_39__N_1404[17] (spi_data_out_r_39__N_1404[17]), 
            .\spi_data_out_r_39__N_1639[17] (spi_data_out_r_39__N_1639[17]), 
            .spi_data_out_r_39__N_6220(spi_data_out_r_39__N_6220), .\spi_data_out_r_39__N_1874[17] (spi_data_out_r_39__N_1874[17]), 
            .\spi_data_out_r_39__N_1169[17] (spi_data_out_r_39__N_1169[17]), 
            .\spi_data_out_r_39__N_2109[17] (spi_data_out_r_39__N_2109[17]), 
            .\spi_data_out_r_39__N_934[17] (spi_data_out_r_39__N_934[17]), 
            .\spi_data_out_r_39__N_2344[17] (spi_data_out_r_39__N_2344[17]), 
            .\spi_data_out_r_39__N_5197[17] (spi_data_out_r_39__N_5197[17]), 
            .\spi_data_out_r_39__N_4854[17] (spi_data_out_r_39__N_4854[17]), 
            .\spi_data_out_r[18] (spi_data_out_r[18]), .\spi_data_out_r_39__N_3825[18] (spi_data_out_r_39__N_3825[18]), 
            .\spi_data_out_r_39__N_4168[18] (spi_data_out_r_39__N_4168[18]), 
            .\spi_data_out_r_39__N_5540[18] (spi_data_out_r_39__N_5540[18]), 
            .\spi_data_out_r_39__N_4511[18] (spi_data_out_r_39__N_4511[18]), 
            .\spi_data_out_r_39__N_1404[18] (spi_data_out_r_39__N_1404[18]), 
            .\spi_data_out_r_39__N_1639[18] (spi_data_out_r_39__N_1639[18]), 
            .\spi_data_out_r_39__N_1874[18] (spi_data_out_r_39__N_1874[18]), 
            .\spi_data_out_r_39__N_1169[18] (spi_data_out_r_39__N_1169[18]), 
            .\spi_data_out_r_39__N_2109[18] (spi_data_out_r_39__N_2109[18]), 
            .\spi_data_out_r_39__N_934[18] (spi_data_out_r_39__N_934[18]), 
            .\spi_data_out_r_39__N_2344[18] (spi_data_out_r_39__N_2344[18]), 
            .\spi_data_out_r_39__N_5197[18] (spi_data_out_r_39__N_5197[18]), 
            .\spi_data_out_r_39__N_4854[18] (spi_data_out_r_39__N_4854[18]), 
            .\spi_data_out_r[19] (spi_data_out_r[19]), .\spi_data_out_r_39__N_3825[19] (spi_data_out_r_39__N_3825[19]), 
            .\spi_data_out_r_39__N_4168[19] (spi_data_out_r_39__N_4168[19]), 
            .\spi_data_out_r_39__N_5540[19] (spi_data_out_r_39__N_5540[19]), 
            .\spi_data_out_r_39__N_4511[19] (spi_data_out_r_39__N_4511[19]), 
            .\spi_data_out_r_39__N_1404[19] (spi_data_out_r_39__N_1404[19]), 
            .\spi_data_out_r_39__N_1639[19] (spi_data_out_r_39__N_1639[19]), 
            .\spi_data_out_r_39__N_1874[19] (spi_data_out_r_39__N_1874[19]), 
            .\spi_data_out_r_39__N_1169[19] (spi_data_out_r_39__N_1169[19]), 
            .\spi_data_out_r_39__N_2109[19] (spi_data_out_r_39__N_2109[19]), 
            .\spi_data_out_r_39__N_934[19] (spi_data_out_r_39__N_934[19]), 
            .\spi_data_out_r_39__N_2344[19] (spi_data_out_r_39__N_2344[19]), 
            .\spi_data_out_r_39__N_5197[19] (spi_data_out_r_39__N_5197[19]), 
            .\spi_data_out_r_39__N_4854[19] (spi_data_out_r_39__N_4854[19]), 
            .\spi_data_out_r[20] (spi_data_out_r[20]), .\spi_data_out_r_39__N_3825[20] (spi_data_out_r_39__N_3825[20]), 
            .\spi_data_out_r_39__N_4168[20] (spi_data_out_r_39__N_4168[20]), 
            .\spi_data_out_r_39__N_5540[20] (spi_data_out_r_39__N_5540[20]), 
            .\spi_data_out_r_39__N_4511[20] (spi_data_out_r_39__N_4511[20]), 
            .\spi_data_out_r_39__N_1404[20] (spi_data_out_r_39__N_1404[20]), 
            .\spi_data_out_r_39__N_1639[20] (spi_data_out_r_39__N_1639[20]), 
            .\spi_data_out_r_39__N_1874[20] (spi_data_out_r_39__N_1874[20]), 
            .\spi_data_out_r_39__N_1169[20] (spi_data_out_r_39__N_1169[20]), 
            .\spi_data_out_r_39__N_2109[20] (spi_data_out_r_39__N_2109[20]), 
            .\spi_data_out_r_39__N_934[20] (spi_data_out_r_39__N_934[20]), 
            .\spi_data_out_r_39__N_2344[20] (spi_data_out_r_39__N_2344[20]), 
            .\spi_data_out_r_39__N_5197[20] (spi_data_out_r_39__N_5197[20]), 
            .\spi_data_out_r_39__N_4854[20] (spi_data_out_r_39__N_4854[20]), 
            .\spi_data_out_r[21] (spi_data_out_r[21]), .\spi_data_out_r_39__N_3825[21] (spi_data_out_r_39__N_3825[21]), 
            .\spi_data_out_r_39__N_4168[21] (spi_data_out_r_39__N_4168[21]), 
            .\spi_data_out_r_39__N_5540[21] (spi_data_out_r_39__N_5540[21]), 
            .\spi_data_out_r_39__N_4511[21] (spi_data_out_r_39__N_4511[21]), 
            .\spi_data_out_r_39__N_1404[21] (spi_data_out_r_39__N_1404[21]), 
            .\spi_data_out_r_39__N_1639[21] (spi_data_out_r_39__N_1639[21]), 
            .\spi_data_out_r_39__N_1874[21] (spi_data_out_r_39__N_1874[21]), 
            .\spi_data_out_r_39__N_1169[21] (spi_data_out_r_39__N_1169[21]), 
            .\spi_data_out_r_39__N_2109[21] (spi_data_out_r_39__N_2109[21]), 
            .\spi_data_out_r_39__N_934[21] (spi_data_out_r_39__N_934[21]), 
            .\spi_data_out_r_39__N_2344[21] (spi_data_out_r_39__N_2344[21]), 
            .\spi_data_out_r_39__N_5197[21] (spi_data_out_r_39__N_5197[21]), 
            .\spi_data_out_r_39__N_4854[21] (spi_data_out_r_39__N_4854[21]), 
            .\spi_data_out_r[22] (spi_data_out_r[22]), .\spi_data_out_r_39__N_3825[22] (spi_data_out_r_39__N_3825[22]), 
            .\spi_data_out_r_39__N_4168[22] (spi_data_out_r_39__N_4168[22]), 
            .\spi_data_out_r_39__N_5540[22] (spi_data_out_r_39__N_5540[22]), 
            .\spi_data_out_r_39__N_4511[22] (spi_data_out_r_39__N_4511[22]), 
            .\spi_data_out_r_39__N_1404[22] (spi_data_out_r_39__N_1404[22]), 
            .\spi_data_out_r_39__N_1639[22] (spi_data_out_r_39__N_1639[22]), 
            .\spi_data_out_r_39__N_1874[22] (spi_data_out_r_39__N_1874[22]), 
            .\spi_data_out_r_39__N_1169[22] (spi_data_out_r_39__N_1169[22]), 
            .\spi_data_out_r_39__N_2109[22] (spi_data_out_r_39__N_2109[22]), 
            .\spi_data_out_r_39__N_934[22] (spi_data_out_r_39__N_934[22]), 
            .\spi_data_out_r_39__N_2344[22] (spi_data_out_r_39__N_2344[22]), 
            .\spi_data_out_r_39__N_5197[22] (spi_data_out_r_39__N_5197[22]), 
            .\spi_data_out_r_39__N_4854[22] (spi_data_out_r_39__N_4854[22]), 
            .\spi_data_out_r[23] (spi_data_out_r[23]), .\spi_data_out_r_39__N_3825[23] (spi_data_out_r_39__N_3825[23]), 
            .\spi_data_out_r_39__N_4168[23] (spi_data_out_r_39__N_4168[23]), 
            .\spi_data_out_r_39__N_5540[23] (spi_data_out_r_39__N_5540[23]), 
            .\spi_data_out_r_39__N_4511[23] (spi_data_out_r_39__N_4511[23]), 
            .\spi_data_out_r_39__N_1404[23] (spi_data_out_r_39__N_1404[23]), 
            .\spi_data_out_r_39__N_1639[23] (spi_data_out_r_39__N_1639[23]), 
            .\spi_data_out_r_39__N_1874[23] (spi_data_out_r_39__N_1874[23]), 
            .\spi_data_out_r_39__N_1169[23] (spi_data_out_r_39__N_1169[23]), 
            .\spi_data_out_r_39__N_2109[23] (spi_data_out_r_39__N_2109[23]), 
            .\spi_data_out_r_39__N_934[23] (spi_data_out_r_39__N_934[23]), 
            .\spi_data_out_r_39__N_2344[23] (spi_data_out_r_39__N_2344[23]), 
            .\spi_data_out_r_39__N_5197[23] (spi_data_out_r_39__N_5197[23]), 
            .\spi_data_out_r_39__N_4854[23] (spi_data_out_r_39__N_4854[23]), 
            .\spi_data_out_r[24] (spi_data_out_r[24]), .\spi_data_out_r_39__N_3825[24] (spi_data_out_r_39__N_3825[24]), 
            .\spi_data_out_r_39__N_4168[24] (spi_data_out_r_39__N_4168[24]), 
            .\spi_data_out_r_39__N_5540[24] (spi_data_out_r_39__N_5540[24]), 
            .\spi_data_out_r_39__N_4511[24] (spi_data_out_r_39__N_4511[24]), 
            .\spi_data_out_r_39__N_1404[24] (spi_data_out_r_39__N_1404[24]), 
            .\spi_data_out_r_39__N_1639[24] (spi_data_out_r_39__N_1639[24]), 
            .\spi_data_out_r_39__N_1874[24] (spi_data_out_r_39__N_1874[24]), 
            .\spi_data_out_r_39__N_1169[24] (spi_data_out_r_39__N_1169[24]), 
            .\spi_data_out_r_39__N_2109[24] (spi_data_out_r_39__N_2109[24]), 
            .\spi_data_out_r_39__N_934[24] (spi_data_out_r_39__N_934[24]), 
            .\spi_data_out_r_39__N_2344[24] (spi_data_out_r_39__N_2344[24]), 
            .\spi_data_out_r_39__N_5197[24] (spi_data_out_r_39__N_5197[24]), 
            .\spi_data_out_r_39__N_4854[24] (spi_data_out_r_39__N_4854[24]), 
            .\spi_data_out_r[25] (spi_data_out_r[25]), .\spi_data_out_r_39__N_3825[25] (spi_data_out_r_39__N_3825[25]), 
            .\spi_data_out_r_39__N_4168[25] (spi_data_out_r_39__N_4168[25]), 
            .\spi_data_out_r_39__N_5540[25] (spi_data_out_r_39__N_5540[25]), 
            .\spi_data_out_r_39__N_4511[25] (spi_data_out_r_39__N_4511[25]), 
            .\spi_data_out_r_39__N_1404[25] (spi_data_out_r_39__N_1404[25]), 
            .\spi_data_out_r_39__N_1639[25] (spi_data_out_r_39__N_1639[25]), 
            .\spi_data_out_r_39__N_1874[25] (spi_data_out_r_39__N_1874[25]), 
            .\spi_data_out_r_39__N_1169[25] (spi_data_out_r_39__N_1169[25]), 
            .\spi_data_out_r_39__N_2109[25] (spi_data_out_r_39__N_2109[25]), 
            .\spi_data_out_r_39__N_934[25] (spi_data_out_r_39__N_934[25]), 
            .\spi_data_out_r_39__N_2344[25] (spi_data_out_r_39__N_2344[25]), 
            .\spi_data_out_r_39__N_5197[25] (spi_data_out_r_39__N_5197[25]), 
            .\spi_data_out_r_39__N_4854[25] (spi_data_out_r_39__N_4854[25]), 
            .\spi_data_out_r[26] (spi_data_out_r[26]), .\spi_data_out_r_39__N_3825[26] (spi_data_out_r_39__N_3825[26]), 
            .\spi_data_out_r_39__N_4168[26] (spi_data_out_r_39__N_4168[26]), 
            .\spi_data_out_r_39__N_5540[26] (spi_data_out_r_39__N_5540[26]), 
            .\spi_data_out_r_39__N_4511[26] (spi_data_out_r_39__N_4511[26]), 
            .\spi_data_out_r_39__N_1404[26] (spi_data_out_r_39__N_1404[26]), 
            .\spi_data_out_r_39__N_1639[26] (spi_data_out_r_39__N_1639[26]), 
            .\spi_data_out_r_39__N_1874[26] (spi_data_out_r_39__N_1874[26]), 
            .\spi_data_out_r_39__N_1169[26] (spi_data_out_r_39__N_1169[26]), 
            .\spi_data_out_r_39__N_2109[26] (spi_data_out_r_39__N_2109[26]), 
            .\spi_data_out_r_39__N_934[26] (spi_data_out_r_39__N_934[26]), 
            .\spi_data_out_r_39__N_2344[26] (spi_data_out_r_39__N_2344[26]), 
            .\spi_data_out_r_39__N_5197[26] (spi_data_out_r_39__N_5197[26]), 
            .\spi_data_out_r_39__N_4854[26] (spi_data_out_r_39__N_4854[26]), 
            .\spi_data_out_r[27] (spi_data_out_r[27]), .\spi_data_out_r_39__N_3825[27] (spi_data_out_r_39__N_3825[27]), 
            .\spi_data_out_r_39__N_4168[27] (spi_data_out_r_39__N_4168[27]), 
            .\spi_data_out_r_39__N_5540[27] (spi_data_out_r_39__N_5540[27]), 
            .\spi_data_out_r_39__N_4511[27] (spi_data_out_r_39__N_4511[27]), 
            .\spi_data_out_r_39__N_1404[27] (spi_data_out_r_39__N_1404[27]), 
            .\spi_data_out_r_39__N_1639[27] (spi_data_out_r_39__N_1639[27]), 
            .\spi_data_out_r_39__N_1874[27] (spi_data_out_r_39__N_1874[27]), 
            .\spi_data_out_r_39__N_1169[27] (spi_data_out_r_39__N_1169[27]), 
            .\spi_data_out_r_39__N_2109[27] (spi_data_out_r_39__N_2109[27]), 
            .\spi_data_out_r_39__N_934[27] (spi_data_out_r_39__N_934[27]), 
            .\spi_data_out_r_39__N_2344[27] (spi_data_out_r_39__N_2344[27]), 
            .\spi_data_out_r_39__N_5197[27] (spi_data_out_r_39__N_5197[27]), 
            .\spi_data_out_r_39__N_4854[27] (spi_data_out_r_39__N_4854[27]), 
            .\spi_data_out_r[28] (spi_data_out_r[28]), .\spi_data_out_r_39__N_3825[28] (spi_data_out_r_39__N_3825[28]), 
            .\spi_data_out_r_39__N_4168[28] (spi_data_out_r_39__N_4168[28]), 
            .\spi_data_out_r_39__N_5540[28] (spi_data_out_r_39__N_5540[28]), 
            .\spi_data_out_r_39__N_4511[28] (spi_data_out_r_39__N_4511[28]), 
            .\spi_data_out_r_39__N_1404[28] (spi_data_out_r_39__N_1404[28]), 
            .\spi_data_out_r_39__N_1639[28] (spi_data_out_r_39__N_1639[28]), 
            .\spi_data_out_r_39__N_1874[28] (spi_data_out_r_39__N_1874[28]), 
            .\spi_data_out_r_39__N_1169[28] (spi_data_out_r_39__N_1169[28]), 
            .\spi_data_out_r_39__N_2109[28] (spi_data_out_r_39__N_2109[28]), 
            .\spi_data_out_r_39__N_934[28] (spi_data_out_r_39__N_934[28]), 
            .\spi_data_out_r_39__N_2344[28] (spi_data_out_r_39__N_2344[28]), 
            .\spi_data_out_r_39__N_5197[28] (spi_data_out_r_39__N_5197[28]), 
            .\spi_data_out_r_39__N_4854[28] (spi_data_out_r_39__N_4854[28]), 
            .\spi_data_out_r[29] (spi_data_out_r[29]), .\spi_data_out_r_39__N_3825[29] (spi_data_out_r_39__N_3825[29]), 
            .\spi_data_out_r_39__N_4168[29] (spi_data_out_r_39__N_4168[29]), 
            .\spi_data_out_r_39__N_5540[29] (spi_data_out_r_39__N_5540[29]), 
            .\spi_data_out_r_39__N_4511[29] (spi_data_out_r_39__N_4511[29]), 
            .\spi_data_out_r_39__N_1404[29] (spi_data_out_r_39__N_1404[29]), 
            .\spi_data_out_r_39__N_1639[29] (spi_data_out_r_39__N_1639[29]), 
            .\spi_data_out_r_39__N_1874[29] (spi_data_out_r_39__N_1874[29]), 
            .\spi_data_out_r_39__N_1169[29] (spi_data_out_r_39__N_1169[29]), 
            .\spi_data_out_r_39__N_2109[29] (spi_data_out_r_39__N_2109[29]), 
            .\spi_data_out_r_39__N_934[29] (spi_data_out_r_39__N_934[29]), 
            .\spi_data_out_r_39__N_2344[29] (spi_data_out_r_39__N_2344[29]), 
            .\spi_data_out_r_39__N_5197[29] (spi_data_out_r_39__N_5197[29]), 
            .\spi_data_out_r_39__N_4854[29] (spi_data_out_r_39__N_4854[29]), 
            .n6(n6), .OW_ID_N_6182(OW_ID_N_6182), .\spi_data_out_r[30] (spi_data_out_r[30]), 
            .\spi_data_out_r_39__N_3825[30] (spi_data_out_r_39__N_3825[30]), 
            .\spi_data_out_r_39__N_4168[30] (spi_data_out_r_39__N_4168[30]), 
            .\spi_data_out_r_39__N_5540[30] (spi_data_out_r_39__N_5540[30]), 
            .\spi_data_out_r_39__N_4511[30] (spi_data_out_r_39__N_4511[30]), 
            .\spi_data_out_r_39__N_1404[30] (spi_data_out_r_39__N_1404[30]), 
            .\spi_data_out_r_39__N_1639[30] (spi_data_out_r_39__N_1639[30]), 
            .\spi_data_out_r_39__N_1874[30] (spi_data_out_r_39__N_1874[30]), 
            .\spi_data_out_r_39__N_1169[30] (spi_data_out_r_39__N_1169[30]), 
            .\spi_data_out_r_39__N_2109[30] (spi_data_out_r_39__N_2109[30]), 
            .\spi_data_out_r_39__N_934[30] (spi_data_out_r_39__N_934[30]), 
            .\spi_data_out_r_39__N_2344[30] (spi_data_out_r_39__N_2344[30]), 
            .\spi_data_out_r_39__N_5197[30] (spi_data_out_r_39__N_5197[30]), 
            .\spi_data_out_r_39__N_4854[30] (spi_data_out_r_39__N_4854[30]), 
            .\spi_data_out_r[31] (spi_data_out_r[31]), .\spi_data_out_r_39__N_3825[31] (spi_data_out_r_39__N_3825[31]), 
            .\spi_data_out_r_39__N_4168[31] (spi_data_out_r_39__N_4168[31]), 
            .\spi_data_out_r_39__N_5540[31] (spi_data_out_r_39__N_5540[31]), 
            .\spi_data_out_r_39__N_4511[31] (spi_data_out_r_39__N_4511[31]), 
            .\spi_data_out_r_39__N_1404[31] (spi_data_out_r_39__N_1404[31]), 
            .\spi_data_out_r_39__N_1639[31] (spi_data_out_r_39__N_1639[31]), 
            .\spi_data_out_r_39__N_1874[31] (spi_data_out_r_39__N_1874[31]), 
            .\spi_data_out_r_39__N_1169[31] (spi_data_out_r_39__N_1169[31]), 
            .\spi_data_out_r_39__N_2109[31] (spi_data_out_r_39__N_2109[31]), 
            .\spi_data_out_r_39__N_934[31] (spi_data_out_r_39__N_934[31]), 
            .\spi_data_out_r_39__N_2344[31] (spi_data_out_r_39__N_2344[31]), 
            .\spi_data_out_r_39__N_5197[31] (spi_data_out_r_39__N_5197[31]), 
            .\spi_data_out_r_39__N_4854[31] (spi_data_out_r_39__N_4854[31]), 
            .\spi_data_out_r_39__N_4168[32] (spi_data_out_r_39__N_4168[32]), 
            .\spi_data_out_r[32] (spi_data_out_r[32]), .\spi_data_out_r_39__N_4854[32] (spi_data_out_r_39__N_4854[32]), 
            .\spi_data_out_r_39__N_5540[32] (spi_data_out_r_39__N_5540[32]), 
            .\spi_data_out_r_39__N_4511[32] (spi_data_out_r_39__N_4511[32]), 
            .\spi_data_out_r_39__N_5197[32] (spi_data_out_r_39__N_5197[32]), 
            .\spi_data_out_r_39__N_3825[32] (spi_data_out_r_39__N_3825[32]), 
            .\spi_data_out_r_39__N_4168[33] (spi_data_out_r_39__N_4168[33]), 
            .\spi_data_out_r[33] (spi_data_out_r[33]), .\spi_data_out_r_39__N_4854[33] (spi_data_out_r_39__N_4854[33]), 
            .\spi_data_out_r_39__N_5540[33] (spi_data_out_r_39__N_5540[33]), 
            .\spi_data_out_r_39__N_4511[33] (spi_data_out_r_39__N_4511[33]), 
            .\spi_data_out_r_39__N_5197[33] (spi_data_out_r_39__N_5197[33]), 
            .\spi_data_out_r_39__N_3825[33] (spi_data_out_r_39__N_3825[33]), 
            .\spi_data_out_r_39__N_4168[34] (spi_data_out_r_39__N_4168[34]), 
            .\spi_data_out_r[34] (spi_data_out_r[34]), .\spi_data_out_r_39__N_4854[34] (spi_data_out_r_39__N_4854[34]), 
            .\spi_data_out_r_39__N_5540[34] (spi_data_out_r_39__N_5540[34]), 
            .\spi_data_out_r_39__N_4511[34] (spi_data_out_r_39__N_4511[34]), 
            .\spi_data_out_r_39__N_5197[34] (spi_data_out_r_39__N_5197[34]), 
            .\spi_data_out_r_39__N_3825[34] (spi_data_out_r_39__N_3825[34]), 
            .\spi_data_out_r_39__N_4168[35] (spi_data_out_r_39__N_4168[35]), 
            .\spi_data_out_r[35] (spi_data_out_r[35]), .\spi_data_out_r_39__N_4854[35] (spi_data_out_r_39__N_4854[35]), 
            .\spi_data_out_r_39__N_5540[35] (spi_data_out_r_39__N_5540[35]), 
            .\spi_data_out_r_39__N_4511[35] (spi_data_out_r_39__N_4511[35]), 
            .\spi_data_out_r_39__N_5197[35] (spi_data_out_r_39__N_5197[35]), 
            .\spi_data_out_r_39__N_3825[35] (spi_data_out_r_39__N_3825[35]), 
            .\spi_data_out_r_39__N_4168[36] (spi_data_out_r_39__N_4168[36]), 
            .\spi_data_out_r[36] (spi_data_out_r[36]), .\spi_data_out_r_39__N_4854[36] (spi_data_out_r_39__N_4854[36]), 
            .\spi_data_out_r_39__N_5540[36] (spi_data_out_r_39__N_5540[36]), 
            .\spi_data_out_r_39__N_4511[36] (spi_data_out_r_39__N_4511[36]), 
            .\spi_data_out_r_39__N_5197[36] (spi_data_out_r_39__N_5197[36]), 
            .\spi_data_out_r_39__N_3825[36] (spi_data_out_r_39__N_3825[36]), 
            .\spi_data_out_r_39__N_4168[37] (spi_data_out_r_39__N_4168[37]), 
            .\spi_data_out_r[37] (spi_data_out_r[37]), .\spi_data_out_r_39__N_4854[37] (spi_data_out_r_39__N_4854[37]), 
            .\spi_data_out_r_39__N_5540[37] (spi_data_out_r_39__N_5540[37]), 
            .\spi_data_out_r_39__N_4511[37] (spi_data_out_r_39__N_4511[37]), 
            .\spi_data_out_r_39__N_5197[37] (spi_data_out_r_39__N_5197[37]), 
            .\spi_data_out_r_39__N_3825[37] (spi_data_out_r_39__N_3825[37]), 
            .\spi_data_out_r_39__N_4168[38] (spi_data_out_r_39__N_4168[38]), 
            .\spi_data_out_r[38] (spi_data_out_r[38]), .\spi_data_out_r_39__N_4854[38] (spi_data_out_r_39__N_4854[38]), 
            .\spi_data_out_r_39__N_5540[38] (spi_data_out_r_39__N_5540[38]), 
            .\spi_data_out_r_39__N_4511[38] (spi_data_out_r_39__N_4511[38]), 
            .\spi_data_out_r_39__N_5197[38] (spi_data_out_r_39__N_5197[38]), 
            .\spi_data_out_r_39__N_3825[38] (spi_data_out_r_39__N_3825[38]), 
            .\spi_data_out_r_39__N_4168[39] (spi_data_out_r_39__N_4168[39]), 
            .\spi_data_out_r[39] (spi_data_out_r[39]), .\spi_data_out_r_39__N_4854[39] (spi_data_out_r_39__N_4854[39]), 
            .\spi_data_out_r_39__N_5540[39] (spi_data_out_r_39__N_5540[39]), 
            .\spi_data_out_r_39__N_4511[39] (spi_data_out_r_39__N_4511[39]), 
            .\spi_data_out_r_39__N_5197[39] (spi_data_out_r_39__N_5197[39]), 
            .\spi_data_out_r_39__N_3825[39] (spi_data_out_r_39__N_3825[39]), 
            .\spi_data_out_r_39__N_5883[8] (spi_data_out_r_39__N_5883[8]), 
            .\spi_data_out_r_39__N_5883[9] (spi_data_out_r_39__N_5883[9]), 
            .n47(n47_adj_7730), .\spi_data_out_r_39__N_3825[8] (spi_data_out_r_39__N_3825[8]), 
            .n16(n16_adj_7461), .\spi_data_out_r_39__N_4511[8] (spi_data_out_r_39__N_4511[8]), 
            .n18(n18_adj_7460), .\spi_data_out_r_39__N_1639[8] (spi_data_out_r_39__N_1639[8]), 
            .n5(n5_adj_7462), .\spi_data_out_r_39__N_1169[8] (spi_data_out_r_39__N_1169[8]), 
            .n3(n3), .\spi_data_out_r_39__N_3825[9] (spi_data_out_r_39__N_3825[9]), 
            .n16_adj_1(n16), .\spi_data_out_r_39__N_5540[9] (spi_data_out_r_39__N_5540[9]), 
            .n21(n21), .\spi_data_out_r_39__N_1639[9] (spi_data_out_r_39__N_1639[9]), 
            .n5_adj_2(n5), .\spi_data_out_r_39__N_934[9] (spi_data_out_r_39__N_934[9]), 
            .n2(n2), .n30165(n30165), .\spi_data_out_r_39__N_5540[2] (spi_data_out_r_39__N_5540[2]), 
            .n21_adj_3(n21_adj_7670), .\spi_data_out_r_39__N_4854[2] (spi_data_out_r_39__N_4854[2]), 
            .n19(n19), .GND_net(GND_net), .\spi_data_out_r_39__N_2109[2] (spi_data_out_r_39__N_2109[2]), 
            .n7(n7), .n22(n22), .\spi_data_out_r_39__N_2934[2] (spi_data_out_r_39__N_2934[2]), 
            .clear_intrpt(clear_intrpt_adj_7665), .n14(n14), .\spi_data_out_r_39__N_2579[2] (spi_data_out_r_39__N_2579[2]), 
            .clear_intrpt_adj_4(clear_intrpt), .n9(n9), .\spi_data_out_r[0] (spi_data_out_r[0]), 
            .\spi_data_out_r_39__N_4854[0] (spi_data_out_r_39__N_4854[0]), 
            .\spi_data_out_r_39__N_4168[0] (spi_data_out_r_39__N_4168[0]), 
            .\spi_data_out_r_39__N_5197[0] (spi_data_out_r_39__N_5197[0]), 
            .\spi_data_out_r_39__N_2650[0] (spi_data_out_r_39__N_2650[0]), 
            .clear_intrpt_adj_5(clear_intrpt_adj_7661), .\spi_data_out_r_39__N_2863[0] (spi_data_out_r_39__N_2863[0]), 
            .clear_intrpt_adj_6(clear_intrpt_adj_7664), .\spi_data_out_r_39__N_2934[0] (spi_data_out_r_39__N_2934[0]), 
            .\spi_data_out_r_39__N_770[0] (spi_data_out_r_39__N_770[0]), .spi_data_out_r_39__N_810(spi_data_out_r_39__N_810), 
            .\spi_data_out_r_39__N_3005[0] (spi_data_out_r_39__N_3005[0]), 
            .clear_intrpt_adj_7(clear_intrpt_adj_7666), .\spi_data_out_r_39__N_2109[0] (spi_data_out_r_39__N_2109[0]), 
            .\spi_data_out_r_39__N_3825[0] (spi_data_out_r_39__N_3825[0]), 
            .\spi_data_out_r_39__N_5540[0] (spi_data_out_r_39__N_5540[0]), 
            .\spi_data_out_r_39__N_2344[0] (spi_data_out_r_39__N_2344[0]), 
            .\spi_data_out_r_39__N_934[0] (spi_data_out_r_39__N_934[0]), .\spi_data_out_r_39__N_1404[0] (spi_data_out_r_39__N_1404[0]), 
            .\spi_data_out_r_39__N_1639[0] (spi_data_out_r_39__N_1639[0]), 
            .\spi_data_out_r_39__N_1169[0] (spi_data_out_r_39__N_1169[0]), 
            .\spi_data_out_r_39__N_1874[0] (spi_data_out_r_39__N_1874[0]), 
            .\spi_data_out_r_39__N_4511[0] (spi_data_out_r_39__N_4511[0]), 
            .\spi_data_out_r_39__N_2792[0] (spi_data_out_r_39__N_2792[0]), 
            .\spi_data_out_r_39__N_2579[0] (spi_data_out_r_39__N_2579[0]), 
            .clear_intrpt_adj_8(clear_intrpt_adj_7663), .\spi_data_out_r_39__N_2721[0] (spi_data_out_r_39__N_2721[0]), 
            .clear_intrpt_adj_9(clear_intrpt_adj_7662), .\uart_slot_en[3] (uart_slot_en[3]), 
            .pin_io_out_65(pin_io_out_65), .n24700(n24700), .pin_io_c_68(pin_io_c_68), 
            .\quad_a[6] (quad_a[6]), .pin_io_out_69(pin_io_out_69), .\quad_b[6] (quad_b[6]), 
            .UC_TXD0_c(UC_TXD0_c), .OW_ID_N_6176(OW_ID_N_6176), .n30083(n30083), 
            .pin_io_c_63(pin_io_c_63), .\pin_intrpt[19] (pin_intrpt[19]), 
            .pin_io_c_64(pin_io_c_64), .\pin_intrpt[20] (pin_intrpt[20]), 
            .pin_io_c_62(pin_io_c_62), .\pin_intrpt[18] (pin_intrpt[18]), 
            .n7258(n7258), .\quad_homing[0] (quad_homing_adj_7967[0]), .n25889(n25889), 
            .\spi_data_out_r[1] (spi_data_out_r[1]), .\spi_data_out_r_39__N_2934[1] (spi_data_out_r_39__N_2934[1]), 
            .\spi_data_out_r_39__N_4511[1] (spi_data_out_r_39__N_4511[1]), 
            .\spi_data_out_r_39__N_5197[1] (spi_data_out_r_39__N_5197[1]), 
            .\spi_data_out_r_39__N_3825[1] (spi_data_out_r_39__N_3825[1]), 
            .\spi_data_out_r_39__N_2863[1] (spi_data_out_r_39__N_2863[1]), 
            .\spi_data_out_r_39__N_3005[1] (spi_data_out_r_39__N_3005[1]), 
            .\spi_data_out_r_39__N_2579[1] (spi_data_out_r_39__N_2579[1]), 
            .\spi_data_out_r_39__N_2792[1] (spi_data_out_r_39__N_2792[1]), 
            .\spi_data_out_r_39__N_2650[1] (spi_data_out_r_39__N_2650[1]), 
            .\spi_data_out_r_39__N_2721[1] (spi_data_out_r_39__N_2721[1]), 
            .\spi_data_out_r_39__N_1169[1] (spi_data_out_r_39__N_1169[1]), 
            .\spi_data_out_r_39__N_4168[1] (spi_data_out_r_39__N_4168[1]), 
            .\spi_data_out_r_39__N_5540[1] (spi_data_out_r_39__N_5540[1]), 
            .\spi_data_out_r_39__N_2344[1] (spi_data_out_r_39__N_2344[1]), 
            .\spi_data_out_r_39__N_1639[1] (spi_data_out_r_39__N_1639[1]), 
            .\spi_data_out_r_39__N_934[1] (spi_data_out_r_39__N_934[1]), .\spi_data_out_r_39__N_2109[1] (spi_data_out_r_39__N_2109[1]), 
            .\spi_data_out_r_39__N_1404[1] (spi_data_out_r_39__N_1404[1]), 
            .\spi_data_out_r_39__N_1874[1] (spi_data_out_r_39__N_1874[1]), 
            .\spi_data_out_r_39__N_4854[1] (spi_data_out_r_39__N_4854[1]), 
            .\spi_data_out_r[3] (spi_data_out_r[3]), .\spi_data_out_r_39__N_3825[3] (spi_data_out_r_39__N_3825[3]), 
            .\spi_data_out_r_39__N_4168[3] (spi_data_out_r_39__N_4168[3]), 
            .\spi_data_out_r_39__N_5540[3] (spi_data_out_r_39__N_5540[3]), 
            .\spi_data_out_r_39__N_4511[3] (spi_data_out_r_39__N_4511[3]), 
            .\spi_data_out_r_39__N_1404[3] (spi_data_out_r_39__N_1404[3]), 
            .\spi_data_out_r_39__N_1639[3] (spi_data_out_r_39__N_1639[3]), 
            .\spi_data_out_r_39__N_1874[3] (spi_data_out_r_39__N_1874[3]), 
            .\spi_data_out_r_39__N_1169[3] (spi_data_out_r_39__N_1169[3]), 
            .\spi_data_out_r_39__N_2109[3] (spi_data_out_r_39__N_2109[3]), 
            .\spi_data_out_r_39__N_934[3] (spi_data_out_r_39__N_934[3]), .\spi_data_out_r_39__N_2344[3] (spi_data_out_r_39__N_2344[3]), 
            .\spi_data_out_r_39__N_5197[3] (spi_data_out_r_39__N_5197[3]), 
            .\spi_data_out_r_39__N_4854[3] (spi_data_out_r_39__N_4854[3]), 
            .\spi_data_out_r[4] (spi_data_out_r[4]), .\spi_data_out_r_39__N_3825[4] (spi_data_out_r_39__N_3825[4]), 
            .\spi_data_out_r_39__N_4168[4] (spi_data_out_r_39__N_4168[4]), 
            .ENC_O_N_6184(ENC_O_N_6184)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(354[3] 397[2])
    \uart_controller(DEV_ID=10,UART_ADDRESS_WIDTH=4)  u_uart_controller (.uart_slot_en({uart_slot_en}), 
            .clk(clk), .clk_enable_320(clk_enable_320), .n30185(n30185), 
            .\spi_data_r[0] (spi_data_r[0]), .spi_cmd_r({spi_cmd_r}), .n23978(n23978), 
            .\spi_data_r[3] (spi_data_r[3]), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[1] (spi_data_r[1]), .\spi_addr_r[3] (spi_addr_r[3]), 
            .spi_data_valid_r(spi_data_valid_r), .\spi_addr_r[0] (spi_addr_r[0]), 
            .n26873(n26873), .\spi_addr_r[1] (spi_addr_r[1]), .n4(n4_adj_7388), 
            .n23916(n23916)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(243[3] 254[2])
    
endmodule
//
// Verilog Description of module \shutter(UART_ADDRESS_WIDTH=4) 
//

module \shutter(UART_ADDRESS_WIDTH=4)  (clk, clk_enable_22, n6590, Phase_4_r, 
            clk_enable_244, n30185, n28546, \spi_cmd_r[3] , n30064, 
            n23916, n26435, clk_enable_695, pwm_duty_2, clk_enable_226, 
            \spi_data_r[0] , n29998, pwm_duty_1, clk_enable_652, pwm_duty_3, 
            clk_enable_738, clk_enable_749, \spi_data_r[11] , \spi_data_r[10] , 
            \spi_data_r[9] , \spi_data_r[8] , \spi_data_r[7] , \spi_data_r[6] , 
            \spi_data_r[5] , Phase_1_r, n28548, \spi_data_r[4] , \spi_data_r[3] , 
            \spi_data_r[2] , \spi_data_r[1] , GND_net, Phase_2_r, n28552, 
            Phase_3_r, n28553, mode, clk_enable_245, clk_enable_613, 
            n6747, \spi_cmd_r[2] , \spi_cmd_r[0] , \spi_addr_r[2] , 
            \spi_addr_r[6] , n26243, \spi_data_r[17] , \spi_data_r[16] , 
            n26521, n21, n19, n20, n26545, \spi_addr_r[4] , n26497, 
            n26569, pwm_out_4_N_6549, pwm_out_1_N_6491, pwm_out_3_N_6530, 
            NSL, n30058, n25347, \pwm_out[0] , mode_adj_660, pwm_out_1, 
            mode_adj_661, reset_r, n30043, n25223, n4, mode_adj_662, 
            digital_output_r, n23148, Phase_r, n24593, UC_TXD0_c, 
            n23409, \uart_slot_en[3] , n30125, \cs_decoded[0] , n11013, 
            n30018, n8, n23722, n23555, n30129, n30052, n24588, 
            pwm_out_2_N_6511, n23610, clk_enable_1105, n6651, clk_enable_1107, 
            n6649, n10500, n7198, n7177, n7201, n30134, n11609, 
            n30175, n11606, n11608, n11008) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input clk_enable_22;
    input n6590;
    output Phase_4_r;
    input clk_enable_244;
    input n30185;
    input n28546;
    input \spi_cmd_r[3] ;
    input n30064;
    input n23916;
    input n26435;
    output clk_enable_695;
    output [11:0]pwm_duty_2;
    input clk_enable_226;
    input \spi_data_r[0] ;
    input n29998;
    output [11:0]pwm_duty_1;
    input clk_enable_652;
    output [11:0]pwm_duty_3;
    input clk_enable_738;
    input clk_enable_749;
    input \spi_data_r[11] ;
    input \spi_data_r[10] ;
    input \spi_data_r[9] ;
    input \spi_data_r[8] ;
    input \spi_data_r[7] ;
    input \spi_data_r[6] ;
    input \spi_data_r[5] ;
    output Phase_1_r;
    input n28548;
    input \spi_data_r[4] ;
    input \spi_data_r[3] ;
    input \spi_data_r[2] ;
    input \spi_data_r[1] ;
    input GND_net;
    output Phase_2_r;
    input n28552;
    output Phase_3_r;
    input n28553;
    output mode;
    input clk_enable_245;
    input clk_enable_613;
    input n6747;
    input \spi_cmd_r[2] ;
    input \spi_cmd_r[0] ;
    input \spi_addr_r[2] ;
    input \spi_addr_r[6] ;
    output n26243;
    input \spi_data_r[17] ;
    input \spi_data_r[16] ;
    output n26521;
    output n21;
    output n19;
    output n20;
    output n26545;
    input \spi_addr_r[4] ;
    output n26497;
    output n26569;
    output pwm_out_4_N_6549;
    output pwm_out_1_N_6491;
    output pwm_out_3_N_6530;
    input NSL;
    input n30058;
    output n25347;
    input \pwm_out[0] ;
    input mode_adj_660;
    input pwm_out_1;
    input mode_adj_661;
    input reset_r;
    input n30043;
    output n25223;
    output n4;
    input [2:0]mode_adj_662;
    input digital_output_r;
    output n23148;
    input Phase_r;
    output n24593;
    input UC_TXD0_c;
    input n23409;
    input \uart_slot_en[3] ;
    output n30125;
    input \cs_decoded[0] ;
    output n11013;
    input n30018;
    input n8;
    input n23722;
    output n23555;
    input n30129;
    input n30052;
    output n24588;
    output pwm_out_2_N_6511;
    output n23610;
    input clk_enable_1105;
    input n6651;
    input clk_enable_1107;
    input n6649;
    output n10500;
    output n7198;
    output n7177;
    output n7201;
    input n30134;
    output n11609;
    input n30175;
    output n11606;
    output n11608;
    output n11008;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    
    wire pwm_out_2;
    wire [11:0]pwm_freq_cntr;   // c:/s_links/sources/slot_cards/shutter_4.v(60[38:51])
    wire [11:0]n53;
    wire [11:0]pwm_duty_4;   // c:/s_links/sources/slot_cards/shutter_4.v(58[38:48])
    
    wire n21912;
    wire [12:0]pwm_out_3_N_6531;
    
    wire n21911, n21986;
    wire [12:0]pwm_out_4_N_6550;
    
    wire n21910, n21985, n21984, n21983, n21982, n21981, n21909, 
        n21790;
    wire [12:0]pwm_out_2_N_6512;
    
    wire n21791, n21908, pwm_out_1_c, n21907, n21801, n21789, n21800, 
        n21788;
    wire [12:0]pwm_out_1_N_6492;
    
    wire n21799, n21798, n21954, n21953, n21787, n21797, n21786, 
        n21796, n21952, n21951, n21950, n21949, n21795, n21794, 
        n21939, n21938, n21937, n21936, n21935, n21934, n6, n3, 
        n30124, n22231, n4_adj_7387, n23740, n25416, n11, n30121, 
        n22225, n21793, n21792, n22132, n22131, n22130, n22129, 
        n22128, pwm_out_3, pwm_out_4, n22127, n28266, n28434, n27107, 
        n28268, n27103;
    
    FD1P3AX pwm_out_2_197 (.D(n6590), .SP(clk_enable_22), .CK(clk), .Q(pwm_out_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(139[8] 199[4])
    defparam pwm_out_2_197.GSR = "DISABLED";
    FD1P3IX Phase_4_r_194 (.D(n28546), .SP(clk_enable_244), .CD(n30185), 
            .CK(clk), .Q(Phase_4_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(115[8] 136[4])
    defparam Phase_4_r_194.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_601_4_lut (.A(\spi_cmd_r[3] ), .B(n30064), .C(n23916), 
         .D(n26435), .Z(clk_enable_695)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_3_lut_rep_601_4_lut.init = 16'h8000;
    FD1P3IX pwm_duty_2__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_226), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_2__i0.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1786__i0 (.D(n53[0]), .CK(clk), .CD(n29998), 
            .Q(pwm_freq_cntr[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786__i0.GSR = "DISABLED";
    FD1P3IX pwm_duty_1__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_652), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_1__i0.GSR = "DISABLED";
    FD1P3IX pwm_duty_3__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_738), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_3[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_3__i0.GSR = "DISABLED";
    FD1P3IX pwm_duty_4__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_749), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_4[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_4__i0.GSR = "DISABLED";
    FD1P3IX pwm_duty_2__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_226), 
            .CD(n30185), .CK(clk), .Q(pwm_duty_2[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_2__i11.GSR = "DISABLED";
    FD1P3IX pwm_duty_2__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_226), 
            .CD(n30185), .CK(clk), .Q(pwm_duty_2[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_2__i10.GSR = "DISABLED";
    FD1P3IX pwm_duty_2__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_226), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_2[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_2__i9.GSR = "DISABLED";
    FD1P3IX pwm_duty_2__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_226), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_2[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_2__i8.GSR = "DISABLED";
    FD1P3IX pwm_duty_2__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_226), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_2[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_2__i7.GSR = "DISABLED";
    FD1P3IX pwm_duty_2__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_226), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_2[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_2__i6.GSR = "DISABLED";
    FD1P3IX pwm_duty_2__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_226), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_2[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_2__i5.GSR = "DISABLED";
    FD1P3IX Phase_1_r_191 (.D(n28548), .SP(clk_enable_244), .CD(n30185), 
            .CK(clk), .Q(Phase_1_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(115[8] 136[4])
    defparam Phase_1_r_191.GSR = "DISABLED";
    FD1P3IX pwm_duty_2__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_226), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_2[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_2__i4.GSR = "DISABLED";
    FD1P3IX pwm_duty_2__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_226), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_2[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_2__i3.GSR = "DISABLED";
    FD1P3IX pwm_duty_2__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_226), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_2__i2.GSR = "DISABLED";
    FD1P3IX pwm_duty_2__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_226), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_2__i1.GSR = "DISABLED";
    CCU2D sub_159_add_2_13 (.A0(pwm_duty_3[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21912), .S0(pwm_out_3_N_6531[11]), .S1(pwm_out_3_N_6531[12]));   // c:/s_links/sources/slot_cards/shutter_4.v(184[25:39])
    defparam sub_159_add_2_13.INIT0 = 16'h5555;
    defparam sub_159_add_2_13.INIT1 = 16'hffff;
    defparam sub_159_add_2_13.INJECT1_0 = "NO";
    defparam sub_159_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_159_add_2_11 (.A0(pwm_duty_3[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_3[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21911), .COUT(n21912), .S0(pwm_out_3_N_6531[9]), 
          .S1(pwm_out_3_N_6531[10]));   // c:/s_links/sources/slot_cards/shutter_4.v(184[25:39])
    defparam sub_159_add_2_11.INIT0 = 16'h5555;
    defparam sub_159_add_2_11.INIT1 = 16'h5555;
    defparam sub_159_add_2_11.INJECT1_0 = "NO";
    defparam sub_159_add_2_11.INJECT1_1 = "NO";
    FD1P3IX Phase_2_r_192 (.D(n28552), .SP(clk_enable_244), .CD(n30185), 
            .CK(clk), .Q(Phase_2_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(115[8] 136[4])
    defparam Phase_2_r_192.GSR = "DISABLED";
    FD1P3IX Phase_3_r_193 (.D(n28553), .SP(clk_enable_244), .CD(n30185), 
            .CK(clk), .Q(Phase_3_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(115[8] 136[4])
    defparam Phase_3_r_193.GSR = "DISABLED";
    FD1P3IX mode_186 (.D(\spi_data_r[0] ), .SP(clk_enable_245), .CD(n30185), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(81[8] 89[4])
    defparam mode_186.GSR = "DISABLED";
    CCU2D sub_164_add_2_13 (.A0(pwm_duty_4[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21986), .S0(pwm_out_4_N_6550[11]), .S1(pwm_out_4_N_6550[12]));   // c:/s_links/sources/slot_cards/shutter_4.v(190[25:39])
    defparam sub_164_add_2_13.INIT0 = 16'h5555;
    defparam sub_164_add_2_13.INIT1 = 16'hffff;
    defparam sub_164_add_2_13.INJECT1_0 = "NO";
    defparam sub_164_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_159_add_2_9 (.A0(pwm_duty_3[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_3[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21910), .COUT(n21911), .S0(pwm_out_3_N_6531[7]), 
          .S1(pwm_out_3_N_6531[8]));   // c:/s_links/sources/slot_cards/shutter_4.v(184[25:39])
    defparam sub_159_add_2_9.INIT0 = 16'h5555;
    defparam sub_159_add_2_9.INIT1 = 16'h5555;
    defparam sub_159_add_2_9.INJECT1_0 = "NO";
    defparam sub_159_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_164_add_2_11 (.A0(pwm_duty_4[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_4[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21985), .COUT(n21986), .S0(pwm_out_4_N_6550[9]), 
          .S1(pwm_out_4_N_6550[10]));   // c:/s_links/sources/slot_cards/shutter_4.v(190[25:39])
    defparam sub_164_add_2_11.INIT0 = 16'h5555;
    defparam sub_164_add_2_11.INIT1 = 16'h5555;
    defparam sub_164_add_2_11.INJECT1_0 = "NO";
    defparam sub_164_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_164_add_2_9 (.A0(pwm_duty_4[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_4[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21984), .COUT(n21985), .S0(pwm_out_4_N_6550[7]), 
          .S1(pwm_out_4_N_6550[8]));   // c:/s_links/sources/slot_cards/shutter_4.v(190[25:39])
    defparam sub_164_add_2_9.INIT0 = 16'h5555;
    defparam sub_164_add_2_9.INIT1 = 16'h5555;
    defparam sub_164_add_2_9.INJECT1_0 = "NO";
    defparam sub_164_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_164_add_2_7 (.A0(pwm_duty_4[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_4[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21983), .COUT(n21984), .S0(pwm_out_4_N_6550[5]), 
          .S1(pwm_out_4_N_6550[6]));   // c:/s_links/sources/slot_cards/shutter_4.v(190[25:39])
    defparam sub_164_add_2_7.INIT0 = 16'h5555;
    defparam sub_164_add_2_7.INIT1 = 16'h5555;
    defparam sub_164_add_2_7.INJECT1_0 = "NO";
    defparam sub_164_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_164_add_2_5 (.A0(pwm_duty_4[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_4[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21982), .COUT(n21983), .S0(pwm_out_4_N_6550[3]), 
          .S1(pwm_out_4_N_6550[4]));   // c:/s_links/sources/slot_cards/shutter_4.v(190[25:39])
    defparam sub_164_add_2_5.INIT0 = 16'h5555;
    defparam sub_164_add_2_5.INIT1 = 16'h5555;
    defparam sub_164_add_2_5.INJECT1_0 = "NO";
    defparam sub_164_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_164_add_2_3 (.A0(pwm_duty_4[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_4[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21981), .COUT(n21982), .S0(pwm_out_4_N_6550[1]), 
          .S1(pwm_out_4_N_6550[2]));   // c:/s_links/sources/slot_cards/shutter_4.v(190[25:39])
    defparam sub_164_add_2_3.INIT0 = 16'h5555;
    defparam sub_164_add_2_3.INIT1 = 16'h5555;
    defparam sub_164_add_2_3.INJECT1_0 = "NO";
    defparam sub_164_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_164_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_duty_4[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n21981), .S1(pwm_out_4_N_6550[0]));   // c:/s_links/sources/slot_cards/shutter_4.v(190[25:39])
    defparam sub_164_add_2_1.INIT0 = 16'hF000;
    defparam sub_164_add_2_1.INIT1 = 16'h5555;
    defparam sub_164_add_2_1.INJECT1_0 = "NO";
    defparam sub_164_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_159_add_2_7 (.A0(pwm_duty_3[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_3[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21909), .COUT(n21910), .S0(pwm_out_3_N_6531[5]), 
          .S1(pwm_out_3_N_6531[6]));   // c:/s_links/sources/slot_cards/shutter_4.v(184[25:39])
    defparam sub_159_add_2_7.INIT0 = 16'h5555;
    defparam sub_159_add_2_7.INIT1 = 16'h5555;
    defparam sub_159_add_2_7.INJECT1_0 = "NO";
    defparam sub_159_add_2_7.INJECT1_1 = "NO";
    CCU2D equal_207_9 (.A0(pwm_out_2_N_6512[11]), .B0(pwm_freq_cntr[11]), 
          .C0(pwm_out_2_N_6512[10]), .D0(pwm_freq_cntr[10]), .A1(pwm_out_2_N_6512[9]), 
          .B1(pwm_freq_cntr[9]), .C1(pwm_out_2_N_6512[8]), .D1(pwm_freq_cntr[8]), 
          .CIN(n21790), .COUT(n21791));
    defparam equal_207_9.INIT0 = 16'h9009;
    defparam equal_207_9.INIT1 = 16'h9009;
    defparam equal_207_9.INJECT1_0 = "YES";
    defparam equal_207_9.INJECT1_1 = "YES";
    CCU2D sub_159_add_2_5 (.A0(pwm_duty_3[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_3[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21908), .COUT(n21909), .S0(pwm_out_3_N_6531[3]), 
          .S1(pwm_out_3_N_6531[4]));   // c:/s_links/sources/slot_cards/shutter_4.v(184[25:39])
    defparam sub_159_add_2_5.INIT0 = 16'h5555;
    defparam sub_159_add_2_5.INIT1 = 16'h5555;
    defparam sub_159_add_2_5.INJECT1_0 = "NO";
    defparam sub_159_add_2_5.INJECT1_1 = "NO";
    CCU2D equal_207_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_out_2_N_6512[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n21790));   // c:/s_links/sources/slot_cards/shutter_4.v(178[8:39])
    defparam equal_207_0.INIT0 = 16'hF000;
    defparam equal_207_0.INIT1 = 16'h5555;
    defparam equal_207_0.INJECT1_0 = "NO";
    defparam equal_207_0.INJECT1_1 = "YES";
    FD1P3AX pwm_out_1_196 (.D(n6747), .SP(clk_enable_613), .CK(clk), .Q(pwm_out_1_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(139[8] 199[4])
    defparam pwm_out_1_196.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1786__i1 (.D(n53[1]), .CK(clk), .CD(n29998), 
            .Q(pwm_freq_cntr[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786__i1.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1786__i2 (.D(n53[2]), .CK(clk), .CD(n29998), 
            .Q(pwm_freq_cntr[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786__i2.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1786__i3 (.D(n53[3]), .CK(clk), .CD(n29998), 
            .Q(pwm_freq_cntr[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786__i3.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1786__i4 (.D(n53[4]), .CK(clk), .CD(n29998), 
            .Q(pwm_freq_cntr[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786__i4.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1786__i5 (.D(n53[5]), .CK(clk), .CD(n29998), 
            .Q(pwm_freq_cntr[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786__i5.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1786__i6 (.D(n53[6]), .CK(clk), .CD(n29998), 
            .Q(pwm_freq_cntr[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786__i6.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1786__i7 (.D(n53[7]), .CK(clk), .CD(n29998), 
            .Q(pwm_freq_cntr[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786__i7.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1786__i8 (.D(n53[8]), .CK(clk), .CD(n29998), 
            .Q(pwm_freq_cntr[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786__i8.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1786__i9 (.D(n53[9]), .CK(clk), .CD(n29998), 
            .Q(pwm_freq_cntr[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786__i9.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1786__i10 (.D(n53[10]), .CK(clk), .CD(n29998), 
            .Q(pwm_freq_cntr[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786__i10.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1786__i11 (.D(n53[11]), .CK(clk), .CD(n29998), 
            .Q(pwm_freq_cntr[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786__i11.GSR = "DISABLED";
    FD1P3IX pwm_duty_1__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_652), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_1__i1.GSR = "DISABLED";
    FD1P3IX pwm_duty_1__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_652), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_1__i2.GSR = "DISABLED";
    FD1P3IX pwm_duty_1__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_652), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_1__i3.GSR = "DISABLED";
    FD1P3IX pwm_duty_1__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_652), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_1__i4.GSR = "DISABLED";
    FD1P3IX pwm_duty_1__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_652), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_1__i5.GSR = "DISABLED";
    FD1P3IX pwm_duty_1__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_652), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_1__i6.GSR = "DISABLED";
    FD1P3IX pwm_duty_1__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_652), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_1__i7.GSR = "DISABLED";
    FD1P3IX pwm_duty_1__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_652), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_1__i8.GSR = "DISABLED";
    FD1P3IX pwm_duty_1__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_652), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_1__i9.GSR = "DISABLED";
    FD1P3IX pwm_duty_1__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_652), 
            .CD(n30185), .CK(clk), .Q(pwm_duty_1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_1__i10.GSR = "DISABLED";
    FD1P3IX pwm_duty_1__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_652), 
            .CD(n30185), .CK(clk), .Q(pwm_duty_1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_1__i11.GSR = "DISABLED";
    CCU2D sub_159_add_2_3 (.A0(pwm_duty_3[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_3[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21907), .COUT(n21908), .S0(pwm_out_3_N_6531[1]), 
          .S1(pwm_out_3_N_6531[2]));   // c:/s_links/sources/slot_cards/shutter_4.v(184[25:39])
    defparam sub_159_add_2_3.INIT0 = 16'h5555;
    defparam sub_159_add_2_3.INIT1 = 16'h5555;
    defparam sub_159_add_2_3.INJECT1_0 = "NO";
    defparam sub_159_add_2_3.INJECT1_1 = "NO";
    FD1P3IX pwm_duty_3__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_738), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_3[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_3__i1.GSR = "DISABLED";
    FD1P3IX pwm_duty_3__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_738), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_3[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_3__i2.GSR = "DISABLED";
    FD1P3IX pwm_duty_3__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_738), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_3[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_3__i3.GSR = "DISABLED";
    FD1P3IX pwm_duty_3__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_738), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_3[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_3__i4.GSR = "DISABLED";
    FD1P3IX pwm_duty_3__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_738), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_3[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_3__i5.GSR = "DISABLED";
    FD1P3IX pwm_duty_3__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_738), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_3[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_3__i6.GSR = "DISABLED";
    FD1P3IX pwm_duty_3__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_738), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_3[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_3__i7.GSR = "DISABLED";
    FD1P3IX pwm_duty_3__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_738), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_3[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_3__i8.GSR = "DISABLED";
    FD1P3IX pwm_duty_3__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_738), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_3[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_3__i9.GSR = "DISABLED";
    FD1P3IX pwm_duty_3__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_738), 
            .CD(n30185), .CK(clk), .Q(pwm_duty_3[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_3__i10.GSR = "DISABLED";
    FD1P3IX pwm_duty_3__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_738), 
            .CD(n30185), .CK(clk), .Q(pwm_duty_3[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_3__i11.GSR = "DISABLED";
    FD1P3IX pwm_duty_4__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_749), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_4[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_4__i1.GSR = "DISABLED";
    FD1P3IX pwm_duty_4__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_749), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_4[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_4__i2.GSR = "DISABLED";
    FD1P3IX pwm_duty_4__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_749), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_4[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_4__i3.GSR = "DISABLED";
    FD1P3IX pwm_duty_4__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_749), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_4[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_4__i4.GSR = "DISABLED";
    FD1P3IX pwm_duty_4__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_749), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_4[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_4__i5.GSR = "DISABLED";
    FD1P3IX pwm_duty_4__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_749), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_4[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_4__i6.GSR = "DISABLED";
    FD1P3IX pwm_duty_4__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_749), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_4[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_4__i7.GSR = "DISABLED";
    FD1P3IX pwm_duty_4__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_749), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_4[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_4__i8.GSR = "DISABLED";
    FD1P3IX pwm_duty_4__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_749), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_4[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_4__i9.GSR = "DISABLED";
    FD1P3IX pwm_duty_4__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_749), 
            .CD(n30185), .CK(clk), .Q(pwm_duty_4[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_4__i10.GSR = "DISABLED";
    FD1P3IX pwm_duty_4__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_749), 
            .CD(n30185), .CK(clk), .Q(pwm_duty_4[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(91[8] 112[4])
    defparam pwm_duty_4__i11.GSR = "DISABLED";
    CCU2D sub_159_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_duty_3[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n21907), .S1(pwm_out_3_N_6531[0]));   // c:/s_links/sources/slot_cards/shutter_4.v(184[25:39])
    defparam sub_159_add_2_1.INIT0 = 16'hF000;
    defparam sub_159_add_2_1.INIT1 = 16'h5555;
    defparam sub_159_add_2_1.INJECT1_0 = "NO";
    defparam sub_159_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut (.A(\spi_cmd_r[2] ), .B(\spi_cmd_r[0] ), .C(\spi_addr_r[2] ), 
         .D(\spi_addr_r[6] ), .Z(n26243)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_3_lut_4_lut_adj_897 (.A(\spi_cmd_r[2] ), .B(\spi_cmd_r[0] ), 
         .C(\spi_data_r[17] ), .D(\spi_data_r[16] ), .Z(n26521)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_897.init = 16'h0080;
    LUT4 i9_4_lut (.A(pwm_duty_4[11]), .B(pwm_duty_4[8]), .C(pwm_duty_4[3]), 
         .D(pwm_duty_4[0]), .Z(n21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(165[8:25])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i7_4_lut (.A(pwm_duty_4[4]), .B(pwm_duty_4[9]), .C(pwm_duty_4[10]), 
         .D(pwm_duty_4[1]), .Z(n19)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(165[8:25])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i8_4_lut (.A(pwm_duty_4[6]), .B(pwm_duty_4[2]), .C(pwm_duty_4[5]), 
         .D(pwm_duty_4[7]), .Z(n20)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(165[8:25])
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut_adj_898 (.A(\spi_cmd_r[2] ), .B(\spi_cmd_r[0] ), 
         .C(\spi_data_r[16] ), .D(\spi_data_r[17] ), .Z(n26545)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_898.init = 16'h0080;
    LUT4 i1_2_lut_3_lut (.A(\spi_cmd_r[2] ), .B(\spi_cmd_r[0] ), .C(\spi_addr_r[4] ), 
         .Z(n26497)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h0808;
    LUT4 i1_3_lut_4_lut_adj_899 (.A(\spi_cmd_r[2] ), .B(\spi_cmd_r[0] ), 
         .C(\spi_data_r[16] ), .D(\spi_data_r[17] ), .Z(n26569)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_899.init = 16'h8000;
    CCU2D equal_209_13 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21801), 
          .S0(pwm_out_4_N_6549));
    defparam equal_209_13.INIT0 = 16'hFFFF;
    defparam equal_209_13.INIT1 = 16'h0000;
    defparam equal_209_13.INJECT1_0 = "NO";
    defparam equal_209_13.INJECT1_1 = "NO";
    CCU2D equal_206_13 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21789), 
          .S0(pwm_out_1_N_6491));
    defparam equal_206_13.INIT0 = 16'hFFFF;
    defparam equal_206_13.INIT1 = 16'h0000;
    defparam equal_206_13.INJECT1_0 = "NO";
    defparam equal_206_13.INJECT1_1 = "NO";
    CCU2D equal_209_13_17471 (.A0(pwm_out_4_N_6550[3]), .B0(pwm_freq_cntr[3]), 
          .C0(pwm_out_4_N_6550[2]), .D0(pwm_freq_cntr[2]), .A1(pwm_out_4_N_6550[1]), 
          .B1(pwm_freq_cntr[1]), .C1(pwm_out_4_N_6550[0]), .D1(pwm_freq_cntr[0]), 
          .CIN(n21800), .COUT(n21801));
    defparam equal_209_13_17471.INIT0 = 16'h9009;
    defparam equal_209_13_17471.INIT1 = 16'h9009;
    defparam equal_209_13_17471.INJECT1_0 = "YES";
    defparam equal_209_13_17471.INJECT1_1 = "YES";
    CCU2D equal_206_13_17468 (.A0(pwm_out_1_N_6492[3]), .B0(pwm_freq_cntr[3]), 
          .C0(pwm_out_1_N_6492[2]), .D0(pwm_freq_cntr[2]), .A1(pwm_out_1_N_6492[1]), 
          .B1(pwm_freq_cntr[1]), .C1(pwm_out_1_N_6492[0]), .D1(pwm_freq_cntr[0]), 
          .CIN(n21788), .COUT(n21789));
    defparam equal_206_13_17468.INIT0 = 16'h9009;
    defparam equal_206_13_17468.INIT1 = 16'h9009;
    defparam equal_206_13_17468.INJECT1_0 = "YES";
    defparam equal_206_13_17468.INJECT1_1 = "YES";
    CCU2D equal_209_11 (.A0(pwm_out_4_N_6550[7]), .B0(pwm_freq_cntr[7]), 
          .C0(pwm_out_4_N_6550[6]), .D0(pwm_freq_cntr[6]), .A1(pwm_out_4_N_6550[5]), 
          .B1(pwm_freq_cntr[5]), .C1(pwm_out_4_N_6550[4]), .D1(pwm_freq_cntr[4]), 
          .CIN(n21799), .COUT(n21800));
    defparam equal_209_11.INIT0 = 16'h9009;
    defparam equal_209_11.INIT1 = 16'h9009;
    defparam equal_209_11.INJECT1_0 = "YES";
    defparam equal_209_11.INJECT1_1 = "YES";
    CCU2D equal_209_9 (.A0(pwm_out_4_N_6550[11]), .B0(pwm_freq_cntr[11]), 
          .C0(pwm_out_4_N_6550[10]), .D0(pwm_freq_cntr[10]), .A1(pwm_out_4_N_6550[9]), 
          .B1(pwm_freq_cntr[9]), .C1(pwm_out_4_N_6550[8]), .D1(pwm_freq_cntr[8]), 
          .CIN(n21798), .COUT(n21799));
    defparam equal_209_9.INIT0 = 16'h9009;
    defparam equal_209_9.INIT1 = 16'h9009;
    defparam equal_209_9.INJECT1_0 = "YES";
    defparam equal_209_9.INJECT1_1 = "YES";
    CCU2D sub_149_add_2_13 (.A0(pwm_duty_1[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21954), .S0(pwm_out_1_N_6492[11]), .S1(pwm_out_1_N_6492[12]));   // c:/s_links/sources/slot_cards/shutter_4.v(172[25:39])
    defparam sub_149_add_2_13.INIT0 = 16'h5555;
    defparam sub_149_add_2_13.INIT1 = 16'hffff;
    defparam sub_149_add_2_13.INJECT1_0 = "NO";
    defparam sub_149_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_149_add_2_11 (.A0(pwm_duty_1[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_1[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21953), .COUT(n21954), .S0(pwm_out_1_N_6492[9]), 
          .S1(pwm_out_1_N_6492[10]));   // c:/s_links/sources/slot_cards/shutter_4.v(172[25:39])
    defparam sub_149_add_2_11.INIT0 = 16'h5555;
    defparam sub_149_add_2_11.INIT1 = 16'h5555;
    defparam sub_149_add_2_11.INJECT1_0 = "NO";
    defparam sub_149_add_2_11.INJECT1_1 = "NO";
    CCU2D equal_209_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_out_4_N_6550[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n21798));   // c:/s_links/sources/slot_cards/shutter_4.v(190[8:39])
    defparam equal_209_0.INIT0 = 16'hF000;
    defparam equal_209_0.INIT1 = 16'h5555;
    defparam equal_209_0.INJECT1_0 = "NO";
    defparam equal_209_0.INJECT1_1 = "YES";
    CCU2D equal_206_11 (.A0(pwm_out_1_N_6492[7]), .B0(pwm_freq_cntr[7]), 
          .C0(pwm_out_1_N_6492[6]), .D0(pwm_freq_cntr[6]), .A1(pwm_out_1_N_6492[5]), 
          .B1(pwm_freq_cntr[5]), .C1(pwm_out_1_N_6492[4]), .D1(pwm_freq_cntr[4]), 
          .CIN(n21787), .COUT(n21788));
    defparam equal_206_11.INIT0 = 16'h9009;
    defparam equal_206_11.INIT1 = 16'h9009;
    defparam equal_206_11.INJECT1_0 = "YES";
    defparam equal_206_11.INJECT1_1 = "YES";
    CCU2D equal_208_13 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21797), 
          .S0(pwm_out_3_N_6530));
    defparam equal_208_13.INIT0 = 16'hFFFF;
    defparam equal_208_13.INIT1 = 16'h0000;
    defparam equal_208_13.INJECT1_0 = "NO";
    defparam equal_208_13.INJECT1_1 = "NO";
    CCU2D equal_206_9 (.A0(pwm_out_1_N_6492[11]), .B0(pwm_freq_cntr[11]), 
          .C0(pwm_out_1_N_6492[10]), .D0(pwm_freq_cntr[10]), .A1(pwm_out_1_N_6492[9]), 
          .B1(pwm_freq_cntr[9]), .C1(pwm_out_1_N_6492[8]), .D1(pwm_freq_cntr[8]), 
          .CIN(n21786), .COUT(n21787));
    defparam equal_206_9.INIT0 = 16'h9009;
    defparam equal_206_9.INIT1 = 16'h9009;
    defparam equal_206_9.INJECT1_0 = "YES";
    defparam equal_206_9.INJECT1_1 = "YES";
    CCU2D equal_208_13_17470 (.A0(pwm_out_3_N_6531[3]), .B0(pwm_freq_cntr[3]), 
          .C0(pwm_out_3_N_6531[2]), .D0(pwm_freq_cntr[2]), .A1(pwm_out_3_N_6531[1]), 
          .B1(pwm_freq_cntr[1]), .C1(pwm_out_3_N_6531[0]), .D1(pwm_freq_cntr[0]), 
          .CIN(n21796), .COUT(n21797));
    defparam equal_208_13_17470.INIT0 = 16'h9009;
    defparam equal_208_13_17470.INIT1 = 16'h9009;
    defparam equal_208_13_17470.INJECT1_0 = "YES";
    defparam equal_208_13_17470.INJECT1_1 = "YES";
    CCU2D equal_206_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_out_1_N_6492[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n21786));   // c:/s_links/sources/slot_cards/shutter_4.v(172[8:39])
    defparam equal_206_0.INIT0 = 16'hF000;
    defparam equal_206_0.INIT1 = 16'h5555;
    defparam equal_206_0.INJECT1_0 = "NO";
    defparam equal_206_0.INJECT1_1 = "YES";
    CCU2D sub_149_add_2_9 (.A0(pwm_duty_1[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_1[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21952), .COUT(n21953), .S0(pwm_out_1_N_6492[7]), 
          .S1(pwm_out_1_N_6492[8]));   // c:/s_links/sources/slot_cards/shutter_4.v(172[25:39])
    defparam sub_149_add_2_9.INIT0 = 16'h5555;
    defparam sub_149_add_2_9.INIT1 = 16'h5555;
    defparam sub_149_add_2_9.INJECT1_0 = "NO";
    defparam sub_149_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_149_add_2_7 (.A0(pwm_duty_1[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_1[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21951), .COUT(n21952), .S0(pwm_out_1_N_6492[5]), 
          .S1(pwm_out_1_N_6492[6]));   // c:/s_links/sources/slot_cards/shutter_4.v(172[25:39])
    defparam sub_149_add_2_7.INIT0 = 16'h5555;
    defparam sub_149_add_2_7.INIT1 = 16'h5555;
    defparam sub_149_add_2_7.INJECT1_0 = "NO";
    defparam sub_149_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_149_add_2_5 (.A0(pwm_duty_1[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_1[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21950), .COUT(n21951), .S0(pwm_out_1_N_6492[3]), 
          .S1(pwm_out_1_N_6492[4]));   // c:/s_links/sources/slot_cards/shutter_4.v(172[25:39])
    defparam sub_149_add_2_5.INIT0 = 16'h5555;
    defparam sub_149_add_2_5.INIT1 = 16'h5555;
    defparam sub_149_add_2_5.INJECT1_0 = "NO";
    defparam sub_149_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_149_add_2_3 (.A0(pwm_duty_1[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_1[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21949), .COUT(n21950), .S0(pwm_out_1_N_6492[1]), 
          .S1(pwm_out_1_N_6492[2]));   // c:/s_links/sources/slot_cards/shutter_4.v(172[25:39])
    defparam sub_149_add_2_3.INIT0 = 16'h5555;
    defparam sub_149_add_2_3.INIT1 = 16'h5555;
    defparam sub_149_add_2_3.INJECT1_0 = "NO";
    defparam sub_149_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_149_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_duty_1[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n21949), .S1(pwm_out_1_N_6492[0]));   // c:/s_links/sources/slot_cards/shutter_4.v(172[25:39])
    defparam sub_149_add_2_1.INIT0 = 16'hF000;
    defparam sub_149_add_2_1.INIT1 = 16'h5555;
    defparam sub_149_add_2_1.INJECT1_0 = "NO";
    defparam sub_149_add_2_1.INJECT1_1 = "NO";
    CCU2D equal_208_11 (.A0(pwm_out_3_N_6531[7]), .B0(pwm_freq_cntr[7]), 
          .C0(pwm_out_3_N_6531[6]), .D0(pwm_freq_cntr[6]), .A1(pwm_out_3_N_6531[5]), 
          .B1(pwm_freq_cntr[5]), .C1(pwm_out_3_N_6531[4]), .D1(pwm_freq_cntr[4]), 
          .CIN(n21795), .COUT(n21796));
    defparam equal_208_11.INIT0 = 16'h9009;
    defparam equal_208_11.INIT1 = 16'h9009;
    defparam equal_208_11.INJECT1_0 = "YES";
    defparam equal_208_11.INJECT1_1 = "YES";
    CCU2D equal_208_9 (.A0(pwm_out_3_N_6531[11]), .B0(pwm_freq_cntr[11]), 
          .C0(pwm_out_3_N_6531[10]), .D0(pwm_freq_cntr[10]), .A1(pwm_out_3_N_6531[9]), 
          .B1(pwm_freq_cntr[9]), .C1(pwm_out_3_N_6531[8]), .D1(pwm_freq_cntr[8]), 
          .CIN(n21794), .COUT(n21795));
    defparam equal_208_9.INIT0 = 16'h9009;
    defparam equal_208_9.INIT1 = 16'h9009;
    defparam equal_208_9.INJECT1_0 = "YES";
    defparam equal_208_9.INJECT1_1 = "YES";
    CCU2D sub_154_add_2_13 (.A0(pwm_duty_2[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21939), .S0(pwm_out_2_N_6512[11]), .S1(pwm_out_2_N_6512[12]));   // c:/s_links/sources/slot_cards/shutter_4.v(178[25:39])
    defparam sub_154_add_2_13.INIT0 = 16'h5555;
    defparam sub_154_add_2_13.INIT1 = 16'hffff;
    defparam sub_154_add_2_13.INJECT1_0 = "NO";
    defparam sub_154_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_154_add_2_11 (.A0(pwm_duty_2[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_2[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21938), .COUT(n21939), .S0(pwm_out_2_N_6512[9]), 
          .S1(pwm_out_2_N_6512[10]));   // c:/s_links/sources/slot_cards/shutter_4.v(178[25:39])
    defparam sub_154_add_2_11.INIT0 = 16'h5555;
    defparam sub_154_add_2_11.INIT1 = 16'h5555;
    defparam sub_154_add_2_11.INJECT1_0 = "NO";
    defparam sub_154_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_154_add_2_9 (.A0(pwm_duty_2[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_2[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21937), .COUT(n21938), .S0(pwm_out_2_N_6512[7]), 
          .S1(pwm_out_2_N_6512[8]));   // c:/s_links/sources/slot_cards/shutter_4.v(178[25:39])
    defparam sub_154_add_2_9.INIT0 = 16'h5555;
    defparam sub_154_add_2_9.INIT1 = 16'h5555;
    defparam sub_154_add_2_9.INJECT1_0 = "NO";
    defparam sub_154_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_154_add_2_7 (.A0(pwm_duty_2[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_2[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21936), .COUT(n21937), .S0(pwm_out_2_N_6512[5]), 
          .S1(pwm_out_2_N_6512[6]));   // c:/s_links/sources/slot_cards/shutter_4.v(178[25:39])
    defparam sub_154_add_2_7.INIT0 = 16'h5555;
    defparam sub_154_add_2_7.INIT1 = 16'h5555;
    defparam sub_154_add_2_7.INJECT1_0 = "NO";
    defparam sub_154_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_154_add_2_5 (.A0(pwm_duty_2[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_2[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21935), .COUT(n21936), .S0(pwm_out_2_N_6512[3]), 
          .S1(pwm_out_2_N_6512[4]));   // c:/s_links/sources/slot_cards/shutter_4.v(178[25:39])
    defparam sub_154_add_2_5.INIT0 = 16'h5555;
    defparam sub_154_add_2_5.INIT1 = 16'h5555;
    defparam sub_154_add_2_5.INJECT1_0 = "NO";
    defparam sub_154_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_154_add_2_3 (.A0(pwm_duty_2[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_2[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21934), .COUT(n21935), .S0(pwm_out_2_N_6512[1]), 
          .S1(pwm_out_2_N_6512[2]));   // c:/s_links/sources/slot_cards/shutter_4.v(178[25:39])
    defparam sub_154_add_2_3.INIT0 = 16'h5555;
    defparam sub_154_add_2_3.INIT1 = 16'h5555;
    defparam sub_154_add_2_3.INJECT1_0 = "NO";
    defparam sub_154_add_2_3.INJECT1_1 = "NO";
    CCU2D equal_208_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_out_3_N_6531[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n21794));   // c:/s_links/sources/slot_cards/shutter_4.v(184[8:39])
    defparam equal_208_0.INIT0 = 16'hF000;
    defparam equal_208_0.INIT1 = 16'h5555;
    defparam equal_208_0.INJECT1_0 = "NO";
    defparam equal_208_0.INJECT1_1 = "YES";
    CCU2D sub_154_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_duty_2[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n21934), .S1(pwm_out_2_N_6512[0]));   // c:/s_links/sources/slot_cards/shutter_4.v(178[25:39])
    defparam sub_154_add_2_1.INIT0 = 16'hF000;
    defparam sub_154_add_2_1.INIT1 = 16'h5555;
    defparam sub_154_add_2_1.INJECT1_0 = "NO";
    defparam sub_154_add_2_1.INJECT1_1 = "NO";
    LUT4 i3_4_lut (.A(NSL), .B(n6), .C(n3), .D(n30058), .Z(n25347)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C))) */ ;
    defparam i3_4_lut.init = 16'hfcfe;
    LUT4 i2_4_lut (.A(Phase_4_r), .B(\pwm_out[0] ), .C(n30124), .D(mode_adj_660), 
         .Z(n6)) /* synthesis lut_function=(A (B (D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i2_4_lut.init = 16'hdc50;
    LUT4 Select_2842_i3_2_lut (.A(pwm_out_1), .B(mode_adj_661), .Z(n3)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2842_i3_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_900 (.A(n22231), .B(mode_adj_661), .C(reset_r), 
         .D(n30043), .Z(n25223)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_900.init = 16'hfeee;
    LUT4 i1_2_lut (.A(mode_adj_660), .B(mode_adj_661), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut (.A(n4_adj_7387), .B(mode_adj_662[1]), .C(n23740), .D(digital_output_r), 
         .Z(n23148)) /* synthesis lut_function=(A+!((C+!(D))+!B)) */ ;
    defparam i1_4_lut.init = 16'haeaa;
    LUT4 Select_2851_i4_2_lut (.A(Phase_r), .B(mode_adj_660), .Z(n4_adj_7387)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2851_i4_2_lut.init = 16'h8888;
    LUT4 i24059_4_lut (.A(n25416), .B(mode_adj_660), .C(mode_adj_662[1]), 
         .D(n23740), .Z(n24593)) /* synthesis lut_function=(!(A+(B+!((D)+!C)))) */ ;
    defparam i24059_4_lut.init = 16'h1101;
    LUT4 i3_4_lut_adj_901 (.A(UC_TXD0_c), .B(n23409), .C(n11), .D(\uart_slot_en[3] ), 
         .Z(n25416)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i3_4_lut_adj_901.init = 16'h0040;
    LUT4 i1_4_lut_adj_902 (.A(n30125), .B(mode_adj_662[2]), .C(mode_adj_662[1]), 
         .D(mode_adj_662[0]), .Z(n11)) /* synthesis lut_function=(!(A (B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_902.init = 16'h5755;
    LUT4 i19116_2_lut (.A(mode_adj_662[2]), .B(mode_adj_662[0]), .Z(n23740)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i19116_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_903 (.A(\cs_decoded[0] ), .B(Phase_3_r), .C(n30043), 
         .D(n30121), .Z(n11013)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_903.init = 16'heca0;
    LUT4 i24062_4_lut (.A(UC_TXD0_c), .B(n30018), .C(n8), .D(n23722), 
         .Z(n23555)) /* synthesis lut_function=(!(A (B)+!A (B+(C (D))))) */ ;
    defparam i24062_4_lut.init = 16'h2333;
    LUT4 i2_4_lut_adj_904 (.A(n22225), .B(mode_adj_661), .C(n30129), .D(n30052), 
         .Z(n24588)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i2_4_lut_adj_904.init = 16'hfeee;
    CCU2D equal_207_13 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21793), 
          .S0(pwm_out_2_N_6511));
    defparam equal_207_13.INIT0 = 16'hFFFF;
    defparam equal_207_13.INIT1 = 16'h0000;
    defparam equal_207_13.INJECT1_0 = "NO";
    defparam equal_207_13.INJECT1_1 = "NO";
    CCU2D equal_207_13_17469 (.A0(pwm_out_2_N_6512[3]), .B0(pwm_freq_cntr[3]), 
          .C0(pwm_out_2_N_6512[2]), .D0(pwm_freq_cntr[2]), .A1(pwm_out_2_N_6512[1]), 
          .B1(pwm_freq_cntr[1]), .C1(pwm_out_2_N_6512[0]), .D1(pwm_freq_cntr[0]), 
          .CIN(n21792), .COUT(n21793));
    defparam equal_207_13_17469.INIT0 = 16'h9009;
    defparam equal_207_13_17469.INIT1 = 16'h9009;
    defparam equal_207_13_17469.INJECT1_0 = "YES";
    defparam equal_207_13_17469.INJECT1_1 = "YES";
    CCU2D equal_207_11 (.A0(pwm_out_2_N_6512[7]), .B0(pwm_freq_cntr[7]), 
          .C0(pwm_out_2_N_6512[6]), .D0(pwm_freq_cntr[6]), .A1(pwm_out_2_N_6512[5]), 
          .B1(pwm_freq_cntr[5]), .C1(pwm_out_2_N_6512[4]), .D1(pwm_freq_cntr[4]), 
          .CIN(n21791), .COUT(n21792));
    defparam equal_207_11.INIT0 = 16'h9009;
    defparam equal_207_11.INIT1 = 16'h9009;
    defparam equal_207_11.INJECT1_0 = "YES";
    defparam equal_207_11.INJECT1_1 = "YES";
    LUT4 i1_3_lut_4_lut_adj_905 (.A(mode_adj_660), .B(n30058), .C(n30125), 
         .D(\cs_decoded[0] ), .Z(n23610)) /* synthesis lut_function=(A+!(B (C+!(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_905.init = 16'hbfbb;
    CCU2D pwm_freq_cntr_1786_add_4_13 (.A0(pwm_freq_cntr[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22132), .S0(n53[11]));   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786_add_4_13.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1786_add_4_13.INIT1 = 16'h0000;
    defparam pwm_freq_cntr_1786_add_4_13.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1786_add_4_13.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1786_add_4_11 (.A0(pwm_freq_cntr[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n22131), .COUT(n22132), .S0(n53[9]), 
          .S1(n53[10]));   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786_add_4_11.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1786_add_4_11.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1786_add_4_11.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1786_add_4_11.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1786_add_4_9 (.A0(pwm_freq_cntr[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n22130), .COUT(n22131), .S0(n53[7]), 
          .S1(n53[8]));   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786_add_4_9.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1786_add_4_9.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1786_add_4_9.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1786_add_4_9.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1786_add_4_7 (.A0(pwm_freq_cntr[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n22129), .COUT(n22130), .S0(n53[5]), 
          .S1(n53[6]));   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786_add_4_7.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1786_add_4_7.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1786_add_4_7.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1786_add_4_7.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1786_add_4_5 (.A0(pwm_freq_cntr[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n22128), .COUT(n22129), .S0(n53[3]), 
          .S1(n53[4]));   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786_add_4_5.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1786_add_4_5.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1786_add_4_5.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1786_add_4_5.INJECT1_1 = "NO";
    FD1P3AX pwm_out_3_198 (.D(n6651), .SP(clk_enable_1105), .CK(clk), 
            .Q(pwm_out_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(139[8] 199[4])
    defparam pwm_out_3_198.GSR = "DISABLED";
    FD1P3AX pwm_out_4_199 (.D(n6649), .SP(clk_enable_1107), .CK(clk), 
            .Q(pwm_out_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=498, LSE_RLINE=530 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(139[8] 199[4])
    defparam pwm_out_4_199.GSR = "DISABLED";
    CCU2D pwm_freq_cntr_1786_add_4_3 (.A0(pwm_freq_cntr[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n22127), .COUT(n22128), .S0(n53[1]), 
          .S1(n53[2]));   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786_add_4_3.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1786_add_4_3.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1786_add_4_3.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1786_add_4_3.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut (.A(mode), .B(pwm_out_2), .C(n4), .D(Phase_2_r), 
         .Z(n10500)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i2_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_3_lut_adj_906 (.A(mode), .B(pwm_out_2), .C(Phase_2_r), 
         .Z(n22225)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_906.init = 16'h0808;
    LUT4 Select_2860_i3_3_lut_4_lut (.A(mode), .B(pwm_out_1_c), .C(Phase_1_r), 
         .D(mode_adj_661), .Z(n7198)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (D)) */ ;
    defparam Select_2860_i3_3_lut_4_lut.init = 16'hff08;
    LUT4 Select_2839_i3_3_lut_4_lut (.A(mode), .B(pwm_out_1_c), .C(mode_adj_661), 
         .D(Phase_1_r), .Z(n7177)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam Select_2839_i3_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i1_2_lut_rep_721 (.A(mode), .B(pwm_out_3), .Z(n30121)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_721.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_907 (.A(mode), .B(pwm_out_3), .C(Phase_3_r), 
         .Z(n22231)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_907.init = 16'h0808;
    LUT4 i1_2_lut_rep_724 (.A(mode), .B(pwm_out_4), .Z(n30124)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_724.init = 16'h8888;
    LUT4 Select_2863_i3_3_lut_4_lut (.A(mode), .B(pwm_out_4), .C(Phase_4_r), 
         .D(mode_adj_661), .Z(n7201)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam Select_2863_i3_3_lut_4_lut.init = 16'hff80;
    LUT4 i24054_2_lut_rep_725 (.A(mode), .B(mode_adj_661), .Z(n30125)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i24054_2_lut_rep_725.init = 16'h1111;
    LUT4 i24045_2_lut_3_lut_4_lut (.A(mode), .B(mode_adj_661), .C(n30134), 
         .D(mode_adj_662[2]), .Z(n11609)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i24045_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i24064_2_lut_3_lut_4_lut (.A(mode), .B(mode_adj_661), .C(mode_adj_662[2]), 
         .D(n30175), .Z(n11606)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i24064_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i24056_2_lut_3_lut (.A(mode), .B(mode_adj_661), .C(mode_adj_660), 
         .Z(n11608)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i24056_2_lut_3_lut.init = 16'h0101;
    CCU2D pwm_freq_cntr_1786_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_freq_cntr[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n22127), .S1(n53[0]));   // c:/s_links/sources/slot_cards/shutter_4.v(196[22:42])
    defparam pwm_freq_cntr_1786_add_4_1.INIT0 = 16'hF000;
    defparam pwm_freq_cntr_1786_add_4_1.INIT1 = 16'h0555;
    defparam pwm_freq_cntr_1786_add_4_1.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1786_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_908 (.A(n28266), .B(n28434), .C(n27107), .D(n28268), 
         .Z(n11008)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i1_4_lut_adj_908.init = 16'hf7ff;
    LUT4 i23564_2_lut (.A(pwm_freq_cntr[5]), .B(pwm_freq_cntr[1]), .Z(n28266)) /* synthesis lut_function=(A (B)) */ ;
    defparam i23564_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_909 (.A(pwm_freq_cntr[3]), .B(pwm_freq_cntr[4]), .C(n27103), 
         .D(pwm_freq_cntr[2]), .Z(n27107)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_909.init = 16'hfffd;
    LUT4 i23566_2_lut (.A(pwm_freq_cntr[0]), .B(pwm_freq_cntr[6]), .Z(n28268)) /* synthesis lut_function=(A (B)) */ ;
    defparam i23566_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_910 (.A(pwm_freq_cntr[11]), .B(pwm_freq_cntr[7]), 
         .Z(n27103)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_910.init = 16'heeee;
    LUT4 i23732_3_lut (.A(pwm_freq_cntr[9]), .B(pwm_freq_cntr[10]), .C(pwm_freq_cntr[8]), 
         .Z(n28434)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i23732_3_lut.init = 16'h8080;
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \intrpt_ctrl(DEV_ID=1) 
//

module \intrpt_ctrl(DEV_ID=1)  (clear_intrpt, clk, n30185, clear_intrpt_N_2717, 
            \spi_data_out_r_39__N_2650[0] , \pin_intrpt[3] , \pin_intrpt[5] , 
            \pin_intrpt[4] , intrpt_out_c_1, intrpt_out_N_2713, n31069, 
            \spi_data_out_r_39__N_2650[2] , \spi_data_out_r_39__N_2650[1] ) /* synthesis syn_module_defined=1 */ ;
    output clear_intrpt;
    input clk;
    input n30185;
    input clear_intrpt_N_2717;
    output \spi_data_out_r_39__N_2650[0] ;
    input \pin_intrpt[3] ;
    input \pin_intrpt[5] ;
    input \pin_intrpt[4] ;
    output intrpt_out_c_1;
    input intrpt_out_N_2713;
    input n31069;
    output \spi_data_out_r_39__N_2650[2] ;
    output \spi_data_out_r_39__N_2650[1] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire \pin_intrpt[5]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[5] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    
    wire assert_intrpt, intrpt_all_edges;
    wire [2:0]intrpt_in_dly;   // c:/s_links/sources/intrpt_ctrl.v(39[36:49])
    wire [2:0]intrpt_in_reg;   // c:/s_links/sources/intrpt_ctrl.v(38[35:48])
    wire [2:0]intrpt_edge;   // c:/s_links/sources/intrpt_ctrl.v(40[36:47])
    
    FD1S3IX clear_intrpt_317 (.D(clear_intrpt_N_2717), .CK(clk), .CD(n30185), 
            .Q(clear_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam clear_intrpt_317.GSR = "DISABLED";
    FD1S3IX assert_intrpt_316 (.D(intrpt_all_edges), .CK(clk), .CD(n30185), 
            .Q(assert_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(63[8] 73[4])
    defparam assert_intrpt_316.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i0 (.D(intrpt_in_reg[0]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\pin_intrpt[3] ), .CK(clk), .Q(\spi_data_out_r_39__N_2650[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i0 (.D(\pin_intrpt[3] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i0.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i2 (.D(\pin_intrpt[5] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i1 (.D(\pin_intrpt[4] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i1.GSR = "DISABLED";
    FD1P3IX intrpt_out_359 (.D(n31069), .SP(assert_intrpt), .CD(intrpt_out_N_2713), 
            .CK(clk), .Q(intrpt_out_c_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(92[8] 99[4])
    defparam intrpt_out_359.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\pin_intrpt[5] ), .CK(clk), .Q(\spi_data_out_r_39__N_2650[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\pin_intrpt[4] ), .CK(clk), .Q(\spi_data_out_r_39__N_2650[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i2 (.D(intrpt_in_reg[2]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i1 (.D(intrpt_in_reg[1]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i1.GSR = "DISABLED";
    LUT4 i2_4_lut (.A(intrpt_edge[2]), .B(intrpt_in_dly[0]), .C(intrpt_edge[1]), 
         .D(intrpt_in_reg[0]), .Z(intrpt_all_edges)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C+(D)))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i2_4_lut.init = 16'hfbfe;
    LUT4 i1400_2_lut (.A(intrpt_in_dly[2]), .B(intrpt_in_reg[2]), .Z(intrpt_edge[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(46[22:89])
    defparam i1400_2_lut.init = 16'h6666;
    LUT4 i1401_2_lut (.A(intrpt_in_dly[1]), .B(intrpt_in_reg[1]), .Z(intrpt_edge[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(46[22:89])
    defparam i1401_2_lut.init = 16'h6666;
    
endmodule
//
// Verilog Description of module \intrpt_ctrl(DEV_ID=2) 
//

module \intrpt_ctrl(DEV_ID=2)  (clk, n30185, \spi_data_out_r_39__N_2721[0] , 
            \pin_intrpt[6] , clear_intrpt, clear_intrpt_N_2788, \pin_intrpt[8] , 
            \pin_intrpt[7] , intrpt_out_c_2, intrpt_out_N_2784, n31069, 
            \spi_data_out_r_39__N_2721[2] , \spi_data_out_r_39__N_2721[1] ) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input n30185;
    output \spi_data_out_r_39__N_2721[0] ;
    input \pin_intrpt[6] ;
    output clear_intrpt;
    input clear_intrpt_N_2788;
    input \pin_intrpt[8] ;
    input \pin_intrpt[7] ;
    output intrpt_out_c_2;
    input intrpt_out_N_2784;
    input n31069;
    output \spi_data_out_r_39__N_2721[2] ;
    output \spi_data_out_r_39__N_2721[1] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire \pin_intrpt[8]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[8] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    wire [2:0]intrpt_in_dly;   // c:/s_links/sources/intrpt_ctrl.v(39[36:49])
    wire [2:0]intrpt_in_reg;   // c:/s_links/sources/intrpt_ctrl.v(38[35:48])
    
    wire assert_intrpt, intrpt_all_edges;
    wire [2:0]intrpt_edge;   // c:/s_links/sources/intrpt_ctrl.v(40[36:47])
    
    FD1S3IX intrpt_in_dly__i0 (.D(intrpt_in_reg[0]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\pin_intrpt[6] ), .CK(clk), .Q(\spi_data_out_r_39__N_2721[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3IX clear_intrpt_317 (.D(clear_intrpt_N_2788), .CK(clk), .CD(n30185), 
            .Q(clear_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam clear_intrpt_317.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i0 (.D(\pin_intrpt[6] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i0.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i2 (.D(\pin_intrpt[8] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i1 (.D(\pin_intrpt[7] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i1.GSR = "DISABLED";
    FD1S3IX assert_intrpt_316 (.D(intrpt_all_edges), .CK(clk), .CD(n30185), 
            .Q(assert_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(63[8] 73[4])
    defparam assert_intrpt_316.GSR = "DISABLED";
    FD1P3IX intrpt_out_359 (.D(n31069), .SP(assert_intrpt), .CD(intrpt_out_N_2784), 
            .CK(clk), .Q(intrpt_out_c_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(92[8] 99[4])
    defparam intrpt_out_359.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\pin_intrpt[8] ), .CK(clk), .Q(\spi_data_out_r_39__N_2721[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\pin_intrpt[7] ), .CK(clk), .Q(\spi_data_out_r_39__N_2721[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i2 (.D(intrpt_in_reg[2]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i1 (.D(intrpt_in_reg[1]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i1.GSR = "DISABLED";
    LUT4 i2_4_lut (.A(intrpt_edge[2]), .B(intrpt_in_dly[0]), .C(intrpt_edge[1]), 
         .D(intrpt_in_reg[0]), .Z(intrpt_all_edges)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C+(D)))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i2_4_lut.init = 16'hfbfe;
    LUT4 i1398_2_lut (.A(intrpt_in_dly[2]), .B(intrpt_in_reg[2]), .Z(intrpt_edge[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(46[22:89])
    defparam i1398_2_lut.init = 16'h6666;
    LUT4 i1399_2_lut (.A(intrpt_in_dly[1]), .B(intrpt_in_reg[1]), .Z(intrpt_edge[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(46[22:89])
    defparam i1399_2_lut.init = 16'h6666;
    
endmodule
//
// Verilog Description of module intrpt_ctrl
//

module intrpt_ctrl (intrpt_out_c_0, clk, intrpt_out_N_2642, n31069, 
            n30185, \spi_data_out_r_39__N_2579[0] , \pin_intrpt[0] , clear_intrpt, 
            \spi_data_out_r_39__N_2579[2] , \pin_intrpt[2] , \spi_data_out_r_39__N_2579[1] , 
            \pin_intrpt[1] , n30198, n30019, n30013, n30027) /* synthesis syn_module_defined=1 */ ;
    output intrpt_out_c_0;
    input clk;
    input intrpt_out_N_2642;
    input n31069;
    input n30185;
    output \spi_data_out_r_39__N_2579[0] ;
    input \pin_intrpt[0] ;
    output clear_intrpt;
    output \spi_data_out_r_39__N_2579[2] ;
    input \pin_intrpt[2] ;
    output \spi_data_out_r_39__N_2579[1] ;
    input \pin_intrpt[1] ;
    input n30198;
    input n30019;
    input n30013;
    input n30027;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire \pin_intrpt[2]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[2] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    
    wire assert_intrpt;
    wire [2:0]intrpt_in_dly;   // c:/s_links/sources/intrpt_ctrl.v(39[36:49])
    wire [2:0]intrpt_in_reg;   // c:/s_links/sources/intrpt_ctrl.v(38[35:48])
    
    wire clear_intrpt_N_2646;
    wire [2:0]intrpt_edge;   // c:/s_links/sources/intrpt_ctrl.v(40[36:47])
    
    wire intrpt_all_edges;
    
    FD1P3IX intrpt_out_359 (.D(n31069), .SP(assert_intrpt), .CD(intrpt_out_N_2642), 
            .CK(clk), .Q(intrpt_out_c_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(92[8] 99[4])
    defparam intrpt_out_359.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i0 (.D(intrpt_in_reg[0]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\pin_intrpt[0] ), .CK(clk), .Q(\spi_data_out_r_39__N_2579[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i0 (.D(\pin_intrpt[0] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i0.GSR = "DISABLED";
    FD1S3IX clear_intrpt_317 (.D(clear_intrpt_N_2646), .CK(clk), .CD(n30185), 
            .Q(clear_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam clear_intrpt_317.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\pin_intrpt[2] ), .CK(clk), .Q(\spi_data_out_r_39__N_2579[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\pin_intrpt[1] ), .CK(clk), .Q(\spi_data_out_r_39__N_2579[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i2 (.D(intrpt_in_reg[2]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i1 (.D(intrpt_in_reg[1]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i1 (.D(\pin_intrpt[1] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i2 (.D(\pin_intrpt[2] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i2.GSR = "DISABLED";
    LUT4 i2_4_lut (.A(intrpt_edge[2]), .B(intrpt_in_dly[0]), .C(intrpt_edge[1]), 
         .D(intrpt_in_reg[0]), .Z(intrpt_all_edges)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C+(D)))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i2_4_lut.init = 16'hfbfe;
    LUT4 i1402_2_lut (.A(intrpt_in_dly[2]), .B(intrpt_in_reg[2]), .Z(intrpt_edge[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(46[22:89])
    defparam i1402_2_lut.init = 16'h6666;
    LUT4 i1404_2_lut (.A(intrpt_in_dly[1]), .B(intrpt_in_reg[1]), .Z(intrpt_edge[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(46[22:89])
    defparam i1404_2_lut.init = 16'h6666;
    LUT4 i24123_4_lut (.A(n30198), .B(n30019), .C(n30013), .D(n30027), 
         .Z(clear_intrpt_N_2646)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(82[15:43])
    defparam i24123_4_lut.init = 16'h0001;
    FD1S3IX assert_intrpt_316 (.D(intrpt_all_edges), .CK(clk), .CD(n30185), 
            .Q(assert_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(63[8] 73[4])
    defparam assert_intrpt_316.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \intrpt_ctrl(DEV_ID=5) 
//

module \intrpt_ctrl(DEV_ID=5)  (clear_intrpt, clk, n30185, clear_intrpt_N_3001, 
            intrpt_out_c_5, intrpt_out_N_2997, n31069, \spi_data_out_r_39__N_2934[0] , 
            \pin_intrpt[15] , \spi_data_out_r_39__N_2934[2] , \pin_intrpt[17] , 
            \spi_data_out_r_39__N_2934[1] , \pin_intrpt[16] ) /* synthesis syn_module_defined=1 */ ;
    output clear_intrpt;
    input clk;
    input n30185;
    input clear_intrpt_N_3001;
    output intrpt_out_c_5;
    input intrpt_out_N_2997;
    input n31069;
    output \spi_data_out_r_39__N_2934[0] ;
    input \pin_intrpt[15] ;
    output \spi_data_out_r_39__N_2934[2] ;
    input \pin_intrpt[17] ;
    output \spi_data_out_r_39__N_2934[1] ;
    input \pin_intrpt[16] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire \pin_intrpt[17]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[17] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    wire [2:0]intrpt_in_dly;   // c:/s_links/sources/intrpt_ctrl.v(39[36:49])
    wire [2:0]intrpt_in_reg;   // c:/s_links/sources/intrpt_ctrl.v(38[35:48])
    wire [2:0]intrpt_edge;   // c:/s_links/sources/intrpt_ctrl.v(40[36:47])
    
    wire assert_intrpt, intrpt_all_edges;
    
    LUT4 i1440_2_lut (.A(intrpt_in_dly[2]), .B(intrpt_in_reg[2]), .Z(intrpt_edge[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(46[22:89])
    defparam i1440_2_lut.init = 16'h6666;
    FD1S3IX clear_intrpt_317 (.D(clear_intrpt_N_3001), .CK(clk), .CD(n30185), 
            .Q(clear_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam clear_intrpt_317.GSR = "DISABLED";
    FD1P3IX intrpt_out_359 (.D(n31069), .SP(assert_intrpt), .CD(intrpt_out_N_2997), 
            .CK(clk), .Q(intrpt_out_c_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(92[8] 99[4])
    defparam intrpt_out_359.GSR = "DISABLED";
    FD1S3IX assert_intrpt_316 (.D(intrpt_all_edges), .CK(clk), .CD(n30185), 
            .Q(assert_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(63[8] 73[4])
    defparam assert_intrpt_316.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i0 (.D(intrpt_in_reg[0]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i0.GSR = "DISABLED";
    LUT4 i1442_2_lut (.A(intrpt_in_dly[1]), .B(intrpt_in_reg[1]), .Z(intrpt_edge[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(46[22:89])
    defparam i1442_2_lut.init = 16'h6666;
    FD1S3AX spi_data_out_r_i1 (.D(\pin_intrpt[15] ), .CK(clk), .Q(\spi_data_out_r_39__N_2934[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i0 (.D(\pin_intrpt[15] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\pin_intrpt[17] ), .CK(clk), .Q(\spi_data_out_r_39__N_2934[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\pin_intrpt[16] ), .CK(clk), .Q(\spi_data_out_r_39__N_2934[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i2 (.D(intrpt_in_reg[2]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i1 (.D(intrpt_in_reg[1]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i1 (.D(\pin_intrpt[16] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i2 (.D(\pin_intrpt[17] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i2.GSR = "DISABLED";
    LUT4 i2_4_lut (.A(intrpt_edge[2]), .B(intrpt_in_dly[0]), .C(intrpt_edge[1]), 
         .D(intrpt_in_reg[0]), .Z(intrpt_all_edges)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C+(D)))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i2_4_lut.init = 16'hfbfe;
    
endmodule
//
// Verilog Description of module \intrpt_ctrl(DEV_ID=3) 
//

module \intrpt_ctrl(DEV_ID=3)  (clk, n30185, \spi_data_out_r_39__N_2792[0] , 
            \pin_intrpt[9] , clear_intrpt, clear_intrpt_N_2859, \pin_intrpt[11] , 
            \pin_intrpt[10] , intrpt_out_c_3, intrpt_out_N_2855, n31069, 
            \spi_data_out_r_39__N_2792[2] , \spi_data_out_r_39__N_2792[1] ) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input n30185;
    output \spi_data_out_r_39__N_2792[0] ;
    input \pin_intrpt[9] ;
    output clear_intrpt;
    input clear_intrpt_N_2859;
    input \pin_intrpt[11] ;
    input \pin_intrpt[10] ;
    output intrpt_out_c_3;
    input intrpt_out_N_2855;
    input n31069;
    output \spi_data_out_r_39__N_2792[2] ;
    output \spi_data_out_r_39__N_2792[1] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire \pin_intrpt[11]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[11] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    wire [2:0]intrpt_in_dly;   // c:/s_links/sources/intrpt_ctrl.v(39[36:49])
    wire [2:0]intrpt_in_reg;   // c:/s_links/sources/intrpt_ctrl.v(38[35:48])
    
    wire assert_intrpt, intrpt_all_edges;
    wire [2:0]intrpt_edge;   // c:/s_links/sources/intrpt_ctrl.v(40[36:47])
    
    FD1S3IX intrpt_in_dly__i0 (.D(intrpt_in_reg[0]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\pin_intrpt[9] ), .CK(clk), .Q(\spi_data_out_r_39__N_2792[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i0 (.D(\pin_intrpt[9] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i0.GSR = "DISABLED";
    FD1S3IX clear_intrpt_317 (.D(clear_intrpt_N_2859), .CK(clk), .CD(n30185), 
            .Q(clear_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam clear_intrpt_317.GSR = "DISABLED";
    FD1S3IX assert_intrpt_316 (.D(intrpt_all_edges), .CK(clk), .CD(n30185), 
            .Q(assert_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(63[8] 73[4])
    defparam assert_intrpt_316.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i2 (.D(\pin_intrpt[11] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i1 (.D(\pin_intrpt[10] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i1.GSR = "DISABLED";
    FD1P3IX intrpt_out_359 (.D(n31069), .SP(assert_intrpt), .CD(intrpt_out_N_2855), 
            .CK(clk), .Q(intrpt_out_c_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(92[8] 99[4])
    defparam intrpt_out_359.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\pin_intrpt[11] ), .CK(clk), .Q(\spi_data_out_r_39__N_2792[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\pin_intrpt[10] ), .CK(clk), .Q(\spi_data_out_r_39__N_2792[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i2 (.D(intrpt_in_reg[2]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i1 (.D(intrpt_in_reg[1]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i1.GSR = "DISABLED";
    LUT4 i2_4_lut (.A(intrpt_edge[2]), .B(intrpt_in_dly[0]), .C(intrpt_edge[1]), 
         .D(intrpt_in_reg[0]), .Z(intrpt_all_edges)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C+(D)))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i2_4_lut.init = 16'hfbfe;
    LUT4 i1396_2_lut (.A(intrpt_in_dly[2]), .B(intrpt_in_reg[2]), .Z(intrpt_edge[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(46[22:89])
    defparam i1396_2_lut.init = 16'h6666;
    LUT4 i1397_2_lut (.A(intrpt_in_dly[1]), .B(intrpt_in_reg[1]), .Z(intrpt_edge[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(46[22:89])
    defparam i1397_2_lut.init = 16'h6666;
    
endmodule
//
// Verilog Description of module cs_decoder
//

module cs_decoder (\cs_decoded[0] , CS_READY_c, n28544, FLASH_CS_c, 
            n30220, MAX3421_CS_c, cs_c_3, cs_c_2, cs_c_4, cs_c_0, 
            cs_c_1, n13, \cs_decoded[12] , n28557, \cs_decoded[10] , 
            n28558, \cs_decoded[8] , n28559, \cs_decoded[6] , n28560, 
            \cs_decoded[4] , n28561, n29575, \cs_decoded_13__N_752[6] , 
            \cs_decoded_13__N_752[0] , n30203, \cs_decoded_13__N_752[10] , 
            n29967, \cs_decoded[2] , n29976, n29977, n30235) /* synthesis syn_module_defined=1 */ ;
    output \cs_decoded[0] ;
    input CS_READY_c;
    input n28544;
    output FLASH_CS_c;
    input n30220;
    output MAX3421_CS_c;
    input cs_c_3;
    input cs_c_2;
    input cs_c_4;
    input cs_c_0;
    input cs_c_1;
    output n13;
    output \cs_decoded[12] ;
    input n28557;
    output \cs_decoded[10] ;
    input n28558;
    output \cs_decoded[8] ;
    input n28559;
    output \cs_decoded[6] ;
    input n28560;
    output \cs_decoded[4] ;
    input n28561;
    output n29575;
    output \cs_decoded_13__N_752[6] ;
    output \cs_decoded_13__N_752[0] ;
    output n30203;
    output \cs_decoded_13__N_752[10] ;
    output n29967;
    output \cs_decoded[2] ;
    output n29976;
    output n29977;
    output n30235;
    
    wire CS_READY_c /* synthesis is_clock=1, SET_AS_NETWORK=CS_READY_c */ ;   // c:/s_links/sources/mcm_top.v(23[24:32])
    
    wire CS_READY_c_enable_8, CS_READY_c_enable_2, CS_READY_c_enable_3, 
        FLASH_CS_N_768, n30119, n30228, n30227, n30231, n30230, 
        n30234, n30233, n29704, CS_READY_c_enable_9;
    wire [13:0]cs_decoded_13__N_752;
    
    FD1P3AY cs_decoded_i0 (.D(n28544), .SP(CS_READY_c_enable_8), .CK(CS_READY_c), 
            .Q(\cs_decoded[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=212 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i0.GSR = "ENABLED";
    FD1P3AY FLASH_CS_14 (.D(n30220), .SP(CS_READY_c_enable_2), .CK(CS_READY_c), 
            .Q(FLASH_CS_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=212 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam FLASH_CS_14.GSR = "ENABLED";
    FD1P3AY MAX3421_CS_15 (.D(FLASH_CS_N_768), .SP(CS_READY_c_enable_3), 
            .CK(CS_READY_c), .Q(MAX3421_CS_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=212 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam MAX3421_CS_15.GSR = "ENABLED";
    LUT4 i24117_2_lut_4_lut (.A(n30119), .B(cs_c_3), .C(cs_c_2), .D(cs_c_4), 
         .Z(CS_READY_c_enable_8)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;   // c:/s_links/sources/cs_decoder.v(32[5] 74[10])
    defparam i24117_2_lut_4_lut.init = 16'h7fff;
    LUT4 i20_3_lut_4_lut_4_lut (.A(cs_c_3), .B(cs_c_0), .C(cs_c_2), .D(cs_c_1), 
         .Z(n13)) /* synthesis lut_function=(A (B (C (D)))+!A (B (C (D))+!B !(C+(D)))) */ ;
    defparam i20_3_lut_4_lut_4_lut.init = 16'hc001;
    FD1P3AY cs_decoded_i12 (.D(n28557), .SP(CS_READY_c_enable_8), .CK(CS_READY_c), 
            .Q(\cs_decoded[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=212 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i12.GSR = "ENABLED";
    FD1P3AY cs_decoded_i10 (.D(n28558), .SP(CS_READY_c_enable_8), .CK(CS_READY_c), 
            .Q(\cs_decoded[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=212 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i10.GSR = "ENABLED";
    FD1P3AY cs_decoded_i8 (.D(n28559), .SP(CS_READY_c_enable_8), .CK(CS_READY_c), 
            .Q(\cs_decoded[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=212 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i8.GSR = "ENABLED";
    FD1P3AY cs_decoded_i6 (.D(n28560), .SP(CS_READY_c_enable_8), .CK(CS_READY_c), 
            .Q(\cs_decoded[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=212 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i6.GSR = "ENABLED";
    FD1P3AY cs_decoded_i4 (.D(n28561), .SP(CS_READY_c_enable_8), .CK(CS_READY_c), 
            .Q(\cs_decoded[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=212 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i4.GSR = "ENABLED";
    LUT4 cs_4__I_0_16_Mux_2_i31_3_lut_then_4_lut (.A(cs_c_4), .B(cs_c_2), 
         .C(cs_c_1), .D(cs_c_3), .Z(n30228)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C (D)+!C !(D))+!B !(C+(D)))) */ ;   // c:/s_links/sources/cs_decoder.v(32[5] 74[10])
    defparam cs_4__I_0_16_Mux_2_i31_3_lut_then_4_lut.init = 16'he2af;
    LUT4 cs_4__I_0_16_Mux_2_i31_3_lut_else_4_lut (.A(cs_c_4), .B(cs_c_2), 
         .C(cs_c_1), .D(cs_c_3), .Z(n30227)) /* synthesis lut_function=(!(A (B (C (D)))+!A (C+(D)))) */ ;   // c:/s_links/sources/cs_decoder.v(32[5] 74[10])
    defparam cs_4__I_0_16_Mux_2_i31_3_lut_else_4_lut.init = 16'h2aaf;
    LUT4 i25_3_lut_then_4_lut (.A(cs_c_4), .B(cs_c_3), .C(cs_c_0), .D(cs_c_1), 
         .Z(n30231)) /* synthesis lut_function=(A ((C (D)+!C !(D))+!B)+!A (B (C (D)))) */ ;
    defparam i25_3_lut_then_4_lut.init = 16'he22a;
    LUT4 i25_3_lut_else_4_lut (.A(cs_c_4), .B(cs_c_3), .C(cs_c_0), .D(cs_c_1), 
         .Z(n30230)) /* synthesis lut_function=(A+!(B+!(C (D)+!C !(D)))) */ ;
    defparam i25_3_lut_else_4_lut.init = 16'hbaab;
    LUT4 i1_4_lut_then_3_lut (.A(cs_c_4), .B(cs_c_0), .C(cs_c_3), .Z(n30234)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i1_4_lut_then_3_lut.init = 16'heaea;
    LUT4 i1_4_lut_else_3_lut (.A(cs_c_4), .B(cs_c_0), .C(cs_c_3), .D(cs_c_1), 
         .Z(n30233)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;
    defparam i1_4_lut_else_3_lut.init = 16'haaab;
    LUT4 cs_c_4_bdd_4_lut (.A(cs_c_4), .B(cs_c_3), .C(cs_c_2), .D(cs_c_1), 
         .Z(n29704)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;
    defparam cs_c_4_bdd_4_lut.init = 16'h8001;
    LUT4 n29704_bdd_2_lut (.A(n29704), .B(cs_c_0), .Z(CS_READY_c_enable_3)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n29704_bdd_2_lut.init = 16'h2222;
    LUT4 i7427_1_lut (.A(cs_c_4), .Z(FLASH_CS_N_768)) /* synthesis lut_function=(!(A)) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i7427_1_lut.init = 16'h5555;
    LUT4 cs_c_1_bdd_4_lut (.A(cs_c_1), .B(cs_c_0), .C(cs_c_3), .D(cs_c_2), 
         .Z(n29575)) /* synthesis lut_function=(A (B (C (D)))+!A !(C+(D))) */ ;
    defparam cs_c_1_bdd_4_lut.init = 16'h8005;
    LUT4 i1_3_lut (.A(cs_c_2), .B(cs_c_4), .C(cs_c_3), .Z(\cs_decoded_13__N_752[6] )) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i1_3_lut.init = 16'hfdfd;
    LUT4 i1_3_lut_adj_896 (.A(cs_c_0), .B(cs_c_4), .C(cs_c_3), .Z(\cs_decoded_13__N_752[0] )) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/s_links/sources/cs_decoder.v(32[5] 74[10])
    defparam i1_3_lut_adj_896.init = 16'hfdfd;
    LUT4 i1_2_lut_rep_803 (.A(cs_c_4), .B(cs_c_3), .Z(n30203)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_803.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut (.A(cs_c_4), .B(cs_c_3), .C(cs_c_2), .Z(\cs_decoded_13__N_752[10] )) /* synthesis lut_function=(A+((C)+!B)) */ ;
    defparam i1_2_lut_3_lut.init = 16'hfbfb;
    LUT4 i4_1_lut (.A(cs_c_1), .Z(CS_READY_c_enable_2)) /* synthesis lut_function=(!(A)) */ ;
    defparam i4_1_lut.init = 16'h5555;
    LUT4 cs_c_3_bdd_4_lut_24389 (.A(cs_c_3), .B(cs_c_1), .C(cs_c_2), .D(cs_c_0), 
         .Z(n29967)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+!(C (D)+!C !(D)))) */ ;
    defparam cs_c_3_bdd_4_lut_24389.init = 16'h9001;
    FD1P3AY cs_decoded_i2 (.D(cs_decoded_13__N_752[2]), .SP(CS_READY_c_enable_9), 
            .CK(CS_READY_c), .Q(\cs_decoded[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=212 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i2.GSR = "ENABLED";
    LUT4 cs_c_3_bdd_4_lut (.A(cs_c_3), .B(cs_c_2), .C(cs_c_0), .D(cs_c_1), 
         .Z(n29976)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A !(B+(C+(D)))) */ ;
    defparam cs_c_3_bdd_4_lut.init = 16'h8021;
    LUT4 i5699_2_lut_rep_719 (.A(cs_c_0), .B(cs_c_1), .Z(n30119)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/cs_decoder.v(32[5] 74[10])
    defparam i5699_2_lut_rep_719.init = 16'h6666;
    LUT4 cs_c_2_bdd_4_lut (.A(cs_c_2), .B(cs_c_0), .C(cs_c_3), .D(cs_c_1), 
         .Z(n29977)) /* synthesis lut_function=(A (B (C (D)))+!A (B (C (D))+!B !(C+(D)))) */ ;
    defparam cs_c_2_bdd_4_lut.init = 16'hc001;
    PFUMX i24403 (.BLUT(n30233), .ALUT(n30234), .C0(cs_c_2), .Z(n30235));
    PFUMX i24401 (.BLUT(n30230), .ALUT(n30231), .C0(cs_c_2), .Z(CS_READY_c_enable_9));
    PFUMX i24399 (.BLUT(n30227), .ALUT(n30228), .C0(cs_c_0), .Z(cs_decoded_13__N_752[2]));
    
endmodule
//
// Verilog Description of module \quad_decoder(DEV_ID=1) 
//

module \quad_decoder(DEV_ID=1)  (quad_homing, clk, clk_enable_520, n30185, 
            \spi_data_r[0] , \quad_a[1] , \quad_b[1] , \spi_data_out_r_39__N_1169[0] , 
            \pin_intrpt[5] , GND_net, clk_enable_842, quad_set_valid_N_1393, 
            spi_data_out_r_39__N_1209, spi_data_out_r_39__N_1398, \spi_data_out_r_39__N_1169[31] , 
            \spi_data_out_r_39__N_1169[30] , \spi_data_out_r_39__N_1169[29] , 
            \spi_data_out_r_39__N_1169[28] , \spi_data_out_r_39__N_1169[27] , 
            \spi_data_out_r_39__N_1169[26] , \spi_data_out_r_39__N_1169[25] , 
            \spi_data_out_r_39__N_1169[24] , \spi_data_out_r_39__N_1169[23] , 
            \spi_data_out_r_39__N_1169[22] , \spi_data_out_r_39__N_1169[21] , 
            \spi_data_out_r_39__N_1169[20] , \spi_data_out_r_39__N_1169[19] , 
            \spi_data_out_r_39__N_1169[18] , \spi_data_out_r_39__N_1169[17] , 
            \spi_data_out_r_39__N_1169[16] , \spi_data_out_r_39__N_1169[15] , 
            \spi_data_out_r_39__N_1169[14] , \spi_data_out_r_39__N_1169[13] , 
            \spi_data_out_r_39__N_1169[12] , \spi_data_out_r_39__N_1169[11] , 
            \spi_data_out_r_39__N_1169[10] , \spi_data_out_r_39__N_1169[9] , 
            \spi_data_out_r_39__N_1169[8] , \spi_data_out_r_39__N_1169[7] , 
            \spi_data_out_r_39__N_1169[6] , \spi_data_out_r_39__N_1169[5] , 
            \spi_data_out_r_39__N_1169[4] , \spi_data_out_r_39__N_1169[3] , 
            \spi_data_out_r_39__N_1169[2] , \spi_data_out_r_39__N_1169[1] , 
            \spi_data_r[1] , n47, \spi_data_r[2] , \spi_data_r[3] , 
            \spi_data_r[4] , \spi_data_r[5] , \spi_data_r[6] , \spi_data_r[7] , 
            \spi_data_r[8] , \spi_data_r[9] , \spi_data_r[10] , \spi_data_r[11] , 
            \spi_data_r[12] , \spi_data_r[13] , \spi_data_r[14] , \spi_data_r[15] , 
            \spi_data_r[16] , \spi_data_r[17] , \spi_data_r[18] , \spi_data_r[19] , 
            \spi_data_r[20] , \spi_data_r[21] , \spi_data_r[22] , \spi_data_r[23] , 
            \spi_data_r[24] , \spi_data_r[25] , \spi_data_r[26] , \spi_data_r[27] , 
            \spi_data_r[28] , \spi_data_r[29] , \spi_data_r[30] , \spi_data_r[31] , 
            n1, resetn_c) /* synthesis syn_module_defined=1 */ ;
    output [1:0]quad_homing;
    input clk;
    input clk_enable_520;
    input n30185;
    input \spi_data_r[0] ;
    input \quad_a[1] ;
    input \quad_b[1] ;
    output \spi_data_out_r_39__N_1169[0] ;
    input \pin_intrpt[5] ;
    input GND_net;
    input clk_enable_842;
    input quad_set_valid_N_1393;
    output spi_data_out_r_39__N_1209;
    input spi_data_out_r_39__N_1398;
    output \spi_data_out_r_39__N_1169[31] ;
    output \spi_data_out_r_39__N_1169[30] ;
    output \spi_data_out_r_39__N_1169[29] ;
    output \spi_data_out_r_39__N_1169[28] ;
    output \spi_data_out_r_39__N_1169[27] ;
    output \spi_data_out_r_39__N_1169[26] ;
    output \spi_data_out_r_39__N_1169[25] ;
    output \spi_data_out_r_39__N_1169[24] ;
    output \spi_data_out_r_39__N_1169[23] ;
    output \spi_data_out_r_39__N_1169[22] ;
    output \spi_data_out_r_39__N_1169[21] ;
    output \spi_data_out_r_39__N_1169[20] ;
    output \spi_data_out_r_39__N_1169[19] ;
    output \spi_data_out_r_39__N_1169[18] ;
    output \spi_data_out_r_39__N_1169[17] ;
    output \spi_data_out_r_39__N_1169[16] ;
    output \spi_data_out_r_39__N_1169[15] ;
    output \spi_data_out_r_39__N_1169[14] ;
    output \spi_data_out_r_39__N_1169[13] ;
    output \spi_data_out_r_39__N_1169[12] ;
    output \spi_data_out_r_39__N_1169[11] ;
    output \spi_data_out_r_39__N_1169[10] ;
    output \spi_data_out_r_39__N_1169[9] ;
    output \spi_data_out_r_39__N_1169[8] ;
    output \spi_data_out_r_39__N_1169[7] ;
    output \spi_data_out_r_39__N_1169[6] ;
    output \spi_data_out_r_39__N_1169[5] ;
    output \spi_data_out_r_39__N_1169[4] ;
    output \spi_data_out_r_39__N_1169[3] ;
    output \spi_data_out_r_39__N_1169[2] ;
    output \spi_data_out_r_39__N_1169[1] ;
    input \spi_data_r[1] ;
    input n47;
    input \spi_data_r[2] ;
    input \spi_data_r[3] ;
    input \spi_data_r[4] ;
    input \spi_data_r[5] ;
    input \spi_data_r[6] ;
    input \spi_data_r[7] ;
    input \spi_data_r[8] ;
    input \spi_data_r[9] ;
    input \spi_data_r[10] ;
    input \spi_data_r[11] ;
    input \spi_data_r[12] ;
    input \spi_data_r[13] ;
    input \spi_data_r[14] ;
    input \spi_data_r[15] ;
    input \spi_data_r[16] ;
    input \spi_data_r[17] ;
    input \spi_data_r[18] ;
    input \spi_data_r[19] ;
    input \spi_data_r[20] ;
    input \spi_data_r[21] ;
    input \spi_data_r[22] ;
    input \spi_data_r[23] ;
    input \spi_data_r[24] ;
    input \spi_data_r[25] ;
    input \spi_data_r[26] ;
    input \spi_data_r[27] ;
    input \spi_data_r[28] ;
    input \spi_data_r[29] ;
    input \spi_data_r[30] ;
    input \spi_data_r[31] ;
    input n1;
    input resetn_c;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire \pin_intrpt[5]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[5] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    wire [31:0]quad_count;   // c:/s_links/sources/quad_decoder.v(43[29:39])
    
    wire clk_enable_519, n8554;
    wire [2:0]quad_a_delayed;   // c:/s_links/sources/quad_decoder.v(34[20:34])
    wire [2:0]quad_b_delayed;   // c:/s_links/sources/quad_decoder.v(35[19:33])
    wire [39:0]spi_data_out_r_39__N_1318;
    wire [31:0]quad_buffer;   // c:/s_links/sources/quad_decoder.v(44[29:40])
    
    wire n22121, n6;
    wire [31:0]n4129;
    
    wire n22122, n22120, n22119, n22118, n22117, n22116, n22115, 
        n22114, n22113, n22112, n22111, n22110, count_dir;
    wire [31:0]quad_set;   // c:/s_links/sources/quad_decoder.v(39[31:39])
    
    wire quad_set_valid, n9821, n9819, n9817, n9815, n9813, n9811, 
        n9809, n9807, n9805, n9803, n9801, n9799, n9797, n9795, 
        n9793, n9791, n9789, n9787, n9785, n9783, n9781, n9779, 
        n9777, n9775, n9773, n9771, n9769, n9767, n9765, n9763, 
        n9761, n5715, n22125, n22124, n22123;
    
    FD1P3IX quad_homing__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_520), .CD(n30185), 
            .CK(clk), .Q(quad_homing[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(62[8] 69[4])
    defparam quad_homing__i0.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i0 (.D(n8554), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i0.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i0 (.D(\quad_a[1] ), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i0.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i0 (.D(\quad_b[1] ), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(spi_data_out_r_39__N_1318[0]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX quad_buffer_i0 (.D(quad_count[0]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i0.GSR = "DISABLED";
    CCU2D add_1361_25 (.A0(quad_count[22]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[23]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22121), .COUT(n22122), .S0(n4129[22]), .S1(n4129[23]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_25.INIT0 = 16'h5569;
    defparam add_1361_25.INIT1 = 16'h5569;
    defparam add_1361_25.INJECT1_0 = "NO";
    defparam add_1361_25.INJECT1_1 = "NO";
    CCU2D add_1361_23 (.A0(quad_count[20]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[21]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22120), .COUT(n22121), .S0(n4129[20]), .S1(n4129[21]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_23.INIT0 = 16'h5569;
    defparam add_1361_23.INIT1 = 16'h5569;
    defparam add_1361_23.INJECT1_0 = "NO";
    defparam add_1361_23.INJECT1_1 = "NO";
    CCU2D add_1361_21 (.A0(quad_count[18]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[19]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22119), .COUT(n22120), .S0(n4129[18]), .S1(n4129[19]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_21.INIT0 = 16'h5569;
    defparam add_1361_21.INIT1 = 16'h5569;
    defparam add_1361_21.INJECT1_0 = "NO";
    defparam add_1361_21.INJECT1_1 = "NO";
    CCU2D add_1361_19 (.A0(quad_count[16]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[17]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22118), .COUT(n22119), .S0(n4129[16]), .S1(n4129[17]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_19.INIT0 = 16'h5569;
    defparam add_1361_19.INIT1 = 16'h5569;
    defparam add_1361_19.INJECT1_0 = "NO";
    defparam add_1361_19.INJECT1_1 = "NO";
    CCU2D add_1361_17 (.A0(quad_count[14]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[15]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22117), .COUT(n22118), .S0(n4129[14]), .S1(n4129[15]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_17.INIT0 = 16'h5569;
    defparam add_1361_17.INIT1 = 16'h5569;
    defparam add_1361_17.INJECT1_0 = "NO";
    defparam add_1361_17.INJECT1_1 = "NO";
    CCU2D add_1361_15 (.A0(quad_count[12]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[13]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22116), .COUT(n22117), .S0(n4129[12]), .S1(n4129[13]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_15.INIT0 = 16'h5569;
    defparam add_1361_15.INIT1 = 16'h5569;
    defparam add_1361_15.INJECT1_0 = "NO";
    defparam add_1361_15.INJECT1_1 = "NO";
    CCU2D add_1361_13 (.A0(quad_count[10]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[11]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22115), .COUT(n22116), .S0(n4129[10]), .S1(n4129[11]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_13.INIT0 = 16'h5569;
    defparam add_1361_13.INIT1 = 16'h5569;
    defparam add_1361_13.INJECT1_0 = "NO";
    defparam add_1361_13.INJECT1_1 = "NO";
    CCU2D add_1361_11 (.A0(quad_count[8]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[9]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22114), .COUT(n22115), .S0(n4129[8]), .S1(n4129[9]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_11.INIT0 = 16'h5569;
    defparam add_1361_11.INIT1 = 16'h5569;
    defparam add_1361_11.INJECT1_0 = "NO";
    defparam add_1361_11.INJECT1_1 = "NO";
    CCU2D add_1361_9 (.A0(quad_count[6]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[7]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22113), .COUT(n22114), .S0(n4129[6]), .S1(n4129[7]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_9.INIT0 = 16'h5569;
    defparam add_1361_9.INIT1 = 16'h5569;
    defparam add_1361_9.INJECT1_0 = "NO";
    defparam add_1361_9.INJECT1_1 = "NO";
    CCU2D add_1361_7 (.A0(quad_count[4]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[5]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22112), .COUT(n22113), .S0(n4129[4]), .S1(n4129[5]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_7.INIT0 = 16'h5569;
    defparam add_1361_7.INIT1 = 16'h5569;
    defparam add_1361_7.INJECT1_0 = "NO";
    defparam add_1361_7.INJECT1_1 = "NO";
    CCU2D add_1361_5 (.A0(quad_count[2]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[3]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22111), .COUT(n22112), .S0(n4129[2]), .S1(n4129[3]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_5.INIT0 = 16'h5569;
    defparam add_1361_5.INIT1 = 16'h5569;
    defparam add_1361_5.INJECT1_0 = "NO";
    defparam add_1361_5.INJECT1_1 = "NO";
    CCU2D add_1361_3 (.A0(quad_count[0]), .B0(count_dir), .C0(n6), .D0(count_dir), 
          .A1(quad_count[1]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22110), .COUT(n22111), .S0(n4129[0]), .S1(n4129[1]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_3.INIT0 = 16'h5665;
    defparam add_1361_3.INIT1 = 16'h5569;
    defparam add_1361_3.INJECT1_0 = "NO";
    defparam add_1361_3.INJECT1_1 = "NO";
    CCU2D add_1361_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quad_a_delayed[2]), .B1(quad_b_delayed[1]), .C1(quad_b_delayed[2]), 
          .D1(quad_a_delayed[1]), .COUT(n22110));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_1.INIT0 = 16'hF000;
    defparam add_1361_1.INIT1 = 16'h0990;
    defparam add_1361_1.INJECT1_0 = "NO";
    defparam add_1361_1.INJECT1_1 = "NO";
    FD1P3IX quad_set__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i0.GSR = "DISABLED";
    FD1S3IX quad_set_valid_388 (.D(quad_set_valid_N_1393), .CK(clk), .CD(n30185), 
            .Q(quad_set_valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set_valid_388.GSR = "DISABLED";
    FD1S3IX i39_391 (.D(spi_data_out_r_39__N_1398), .CK(clk), .CD(n30185), 
            .Q(spi_data_out_r_39__N_1209)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam i39_391.GSR = "DISABLED";
    FD1S3AX quad_buffer_i31 (.D(quad_count[31]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i31.GSR = "DISABLED";
    FD1S3AX quad_buffer_i30 (.D(quad_count[30]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i30.GSR = "DISABLED";
    FD1S3AX quad_buffer_i29 (.D(quad_count[29]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i29.GSR = "DISABLED";
    FD1S3AX quad_buffer_i28 (.D(quad_count[28]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i28.GSR = "DISABLED";
    FD1S3AX quad_buffer_i27 (.D(quad_count[27]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i27.GSR = "DISABLED";
    FD1S3AX quad_buffer_i26 (.D(quad_count[26]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i26.GSR = "DISABLED";
    FD1S3AX quad_buffer_i25 (.D(quad_count[25]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i25.GSR = "DISABLED";
    FD1S3AX quad_buffer_i24 (.D(quad_count[24]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i24.GSR = "DISABLED";
    FD1S3AX quad_buffer_i23 (.D(quad_count[23]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i23.GSR = "DISABLED";
    FD1S3AX quad_buffer_i22 (.D(quad_count[22]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i22.GSR = "DISABLED";
    FD1S3AX quad_buffer_i21 (.D(quad_count[21]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i21.GSR = "DISABLED";
    FD1S3AX quad_buffer_i20 (.D(quad_count[20]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i20.GSR = "DISABLED";
    FD1S3AX quad_buffer_i19 (.D(quad_count[19]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i19.GSR = "DISABLED";
    FD1S3AX quad_buffer_i18 (.D(quad_count[18]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i18.GSR = "DISABLED";
    FD1S3AX quad_buffer_i17 (.D(quad_count[17]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i17.GSR = "DISABLED";
    FD1S3AX quad_buffer_i16 (.D(quad_count[16]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i16.GSR = "DISABLED";
    FD1S3AX quad_buffer_i15 (.D(quad_count[15]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i15.GSR = "DISABLED";
    FD1S3AX quad_buffer_i14 (.D(quad_count[14]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i14.GSR = "DISABLED";
    FD1S3AX quad_buffer_i13 (.D(quad_count[13]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i13.GSR = "DISABLED";
    FD1S3AX quad_buffer_i12 (.D(quad_count[12]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i12.GSR = "DISABLED";
    FD1S3AX quad_buffer_i11 (.D(quad_count[11]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i11.GSR = "DISABLED";
    FD1S3AX quad_buffer_i10 (.D(quad_count[10]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i10.GSR = "DISABLED";
    FD1S3AX quad_buffer_i9 (.D(quad_count[9]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i9.GSR = "DISABLED";
    FD1S3AX quad_buffer_i8 (.D(quad_count[8]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i8.GSR = "DISABLED";
    FD1S3AX quad_buffer_i7 (.D(quad_count[7]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i7.GSR = "DISABLED";
    FD1S3AX quad_buffer_i6 (.D(quad_count[6]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i6.GSR = "DISABLED";
    FD1S3AX quad_buffer_i5 (.D(quad_count[5]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i5.GSR = "DISABLED";
    FD1S3AX quad_buffer_i4 (.D(quad_count[4]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i4.GSR = "DISABLED";
    FD1S3AX quad_buffer_i3 (.D(quad_count[3]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i3.GSR = "DISABLED";
    FD1S3AX quad_buffer_i2 (.D(quad_count[2]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i2.GSR = "DISABLED";
    FD1S3AX quad_buffer_i1 (.D(quad_count[1]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(spi_data_out_r_39__N_1318[31]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i31 (.D(spi_data_out_r_39__N_1318[30]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i30 (.D(spi_data_out_r_39__N_1318[29]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i29 (.D(spi_data_out_r_39__N_1318[28]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i28 (.D(spi_data_out_r_39__N_1318[27]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i27 (.D(spi_data_out_r_39__N_1318[26]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i26 (.D(spi_data_out_r_39__N_1318[25]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i25 (.D(spi_data_out_r_39__N_1318[24]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i24 (.D(spi_data_out_r_39__N_1318[23]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i23 (.D(spi_data_out_r_39__N_1318[22]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i22 (.D(spi_data_out_r_39__N_1318[21]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i21 (.D(spi_data_out_r_39__N_1318[20]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i20 (.D(spi_data_out_r_39__N_1318[19]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i19 (.D(spi_data_out_r_39__N_1318[18]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i18 (.D(spi_data_out_r_39__N_1318[17]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i17 (.D(spi_data_out_r_39__N_1318[16]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i16 (.D(spi_data_out_r_39__N_1318[15]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(spi_data_out_r_39__N_1318[14]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(spi_data_out_r_39__N_1318[13]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(spi_data_out_r_39__N_1318[12]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(spi_data_out_r_39__N_1318[11]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(spi_data_out_r_39__N_1318[10]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(spi_data_out_r_39__N_1318[9]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(spi_data_out_r_39__N_1318[8]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(spi_data_out_r_39__N_1318[7]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(spi_data_out_r_39__N_1318[6]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(spi_data_out_r_39__N_1318[5]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(spi_data_out_r_39__N_1318[4]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(spi_data_out_r_39__N_1318[3]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(spi_data_out_r_39__N_1318[2]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(spi_data_out_r_39__N_1318[1]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1169[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i2 (.D(quad_b_delayed[1]), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i2.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i1 (.D(quad_b_delayed[0]), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i1.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i2 (.D(quad_a_delayed[1]), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i2.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i1 (.D(quad_a_delayed[0]), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i1.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i31 (.D(n9821), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i31.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i30 (.D(n9819), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i30.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i29 (.D(n9817), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i29.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i28 (.D(n9815), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i28.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i27 (.D(n9813), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i27.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i26 (.D(n9811), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i26.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i25 (.D(n9809), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i25.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i24 (.D(n9807), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i24.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i23 (.D(n9805), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i23.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i22 (.D(n9803), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i22.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i21 (.D(n9801), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i21.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i20 (.D(n9799), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i20.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i19 (.D(n9797), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i19.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i18 (.D(n9795), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i18.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i17 (.D(n9793), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i17.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i16 (.D(n9791), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i16.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i15 (.D(n9789), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i15.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i14 (.D(n9787), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i14.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i13 (.D(n9785), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i13.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i12 (.D(n9783), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i12.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i11 (.D(n9781), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i11.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i10 (.D(n9779), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i10.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i9 (.D(n9777), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i9.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i8 (.D(n9775), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i8.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i7 (.D(n9773), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i7.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i6 (.D(n9771), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i6.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i5 (.D(n9769), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i5.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i4 (.D(n9767), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i4.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i3 (.D(n9765), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i3.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i2 (.D(n9763), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i1 (.D(n9761), .SP(clk_enable_519), .CK(clk), 
            .Q(quad_count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i1.GSR = "DISABLED";
    FD1P3IX quad_homing__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_520), .CD(n30185), 
            .CK(clk), .Q(quad_homing[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(62[8] 69[4])
    defparam quad_homing__i1.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(quad_a_delayed[1]), .B(quad_b_delayed[2]), .Z(count_dir)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(96[19:96])
    defparam i1_2_lut.init = 16'h6666;
    LUT4 mux_423_i1_3_lut (.A(quad_count[0]), .B(quad_buffer[0]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i1_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut (.A(quad_b_delayed[1]), .B(quad_a_delayed[2]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(96[19:96])
    defparam i2_2_lut.init = 16'h6666;
    LUT4 mux_423_i32_3_lut (.A(quad_count[31]), .B(quad_buffer[31]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i32_3_lut.init = 16'hcaca;
    LUT4 mux_423_i31_3_lut (.A(quad_count[30]), .B(quad_buffer[30]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i31_3_lut.init = 16'hcaca;
    LUT4 mux_423_i30_3_lut (.A(quad_count[29]), .B(quad_buffer[29]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i30_3_lut.init = 16'hcaca;
    LUT4 mux_423_i29_3_lut (.A(quad_count[28]), .B(quad_buffer[28]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i29_3_lut.init = 16'hcaca;
    LUT4 mux_423_i28_3_lut (.A(quad_count[27]), .B(quad_buffer[27]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i28_3_lut.init = 16'hcaca;
    LUT4 mux_423_i27_3_lut (.A(quad_count[26]), .B(quad_buffer[26]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i27_3_lut.init = 16'hcaca;
    FD1P3IX quad_set__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i1.GSR = "DISABLED";
    FD1P3IX quad_set__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i2.GSR = "DISABLED";
    FD1P3IX quad_set__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i3.GSR = "DISABLED";
    FD1P3IX quad_set__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i4.GSR = "DISABLED";
    FD1P3IX quad_set__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i5.GSR = "DISABLED";
    FD1P3IX quad_set__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i6.GSR = "DISABLED";
    FD1P3IX quad_set__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i7.GSR = "DISABLED";
    FD1P3IX quad_set__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i8.GSR = "DISABLED";
    FD1P3IX quad_set__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i9.GSR = "DISABLED";
    FD1P3IX quad_set__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i10.GSR = "DISABLED";
    FD1P3IX quad_set__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i11.GSR = "DISABLED";
    FD1P3IX quad_set__i12 (.D(\spi_data_r[12] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i12.GSR = "DISABLED";
    FD1P3IX quad_set__i13 (.D(\spi_data_r[13] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i13.GSR = "DISABLED";
    FD1P3IX quad_set__i14 (.D(\spi_data_r[14] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i14.GSR = "DISABLED";
    FD1P3IX quad_set__i15 (.D(\spi_data_r[15] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i15.GSR = "DISABLED";
    FD1P3IX quad_set__i16 (.D(\spi_data_r[16] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i16.GSR = "DISABLED";
    FD1P3IX quad_set__i17 (.D(\spi_data_r[17] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i17.GSR = "DISABLED";
    FD1P3IX quad_set__i18 (.D(\spi_data_r[18] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i18.GSR = "DISABLED";
    FD1P3IX quad_set__i19 (.D(\spi_data_r[19] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i19.GSR = "DISABLED";
    FD1P3IX quad_set__i20 (.D(\spi_data_r[20] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i20.GSR = "DISABLED";
    FD1P3IX quad_set__i21 (.D(\spi_data_r[21] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i21.GSR = "DISABLED";
    FD1P3IX quad_set__i22 (.D(\spi_data_r[22] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i22.GSR = "DISABLED";
    FD1P3IX quad_set__i23 (.D(\spi_data_r[23] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i23.GSR = "DISABLED";
    FD1P3IX quad_set__i24 (.D(\spi_data_r[24] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i24.GSR = "DISABLED";
    FD1P3IX quad_set__i25 (.D(\spi_data_r[25] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i25.GSR = "DISABLED";
    FD1P3IX quad_set__i26 (.D(\spi_data_r[26] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i26.GSR = "DISABLED";
    FD1P3IX quad_set__i27 (.D(\spi_data_r[27] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i27.GSR = "DISABLED";
    FD1P3IX quad_set__i28 (.D(\spi_data_r[28] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i28.GSR = "DISABLED";
    FD1P3IX quad_set__i29 (.D(\spi_data_r[29] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i29.GSR = "DISABLED";
    FD1P3IX quad_set__i30 (.D(\spi_data_r[30] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i30.GSR = "DISABLED";
    FD1P3IX quad_set__i31 (.D(\spi_data_r[31] ), .SP(clk_enable_842), .CD(n30185), 
            .CK(clk), .Q(quad_set[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i31.GSR = "DISABLED";
    LUT4 mux_423_i26_3_lut (.A(quad_count[25]), .B(quad_buffer[25]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i26_3_lut.init = 16'hcaca;
    LUT4 mux_423_i25_3_lut (.A(quad_count[24]), .B(quad_buffer[24]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i25_3_lut.init = 16'hcaca;
    LUT4 mux_423_i24_3_lut (.A(quad_count[23]), .B(quad_buffer[23]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i24_3_lut.init = 16'hcaca;
    LUT4 mux_423_i23_3_lut (.A(quad_count[22]), .B(quad_buffer[22]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i23_3_lut.init = 16'hcaca;
    LUT4 mux_423_i22_3_lut (.A(quad_count[21]), .B(quad_buffer[21]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i22_3_lut.init = 16'hcaca;
    LUT4 mux_423_i21_3_lut (.A(quad_count[20]), .B(quad_buffer[20]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i21_3_lut.init = 16'hcaca;
    LUT4 mux_423_i20_3_lut (.A(quad_count[19]), .B(quad_buffer[19]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i20_3_lut.init = 16'hcaca;
    LUT4 mux_423_i19_3_lut (.A(quad_count[18]), .B(quad_buffer[18]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i19_3_lut.init = 16'hcaca;
    LUT4 mux_423_i18_3_lut (.A(quad_count[17]), .B(quad_buffer[17]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i18_3_lut.init = 16'hcaca;
    LUT4 mux_423_i17_3_lut (.A(quad_count[16]), .B(quad_buffer[16]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i17_3_lut.init = 16'hcaca;
    LUT4 mux_423_i16_3_lut (.A(quad_count[15]), .B(quad_buffer[15]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i16_3_lut.init = 16'hcaca;
    LUT4 mux_423_i15_3_lut (.A(quad_count[14]), .B(quad_buffer[14]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i15_3_lut.init = 16'hcaca;
    LUT4 i4230_4_lut (.A(n4129[0]), .B(quad_set[0]), .C(n5715), .D(n1), 
         .Z(n8554)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4230_4_lut.init = 16'hc0ca;
    LUT4 mux_423_i14_3_lut (.A(quad_count[13]), .B(quad_buffer[13]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i14_3_lut.init = 16'hcaca;
    LUT4 mux_423_i13_3_lut (.A(quad_count[12]), .B(quad_buffer[12]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i13_3_lut.init = 16'hcaca;
    LUT4 mux_423_i12_3_lut (.A(quad_count[11]), .B(quad_buffer[11]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i12_3_lut.init = 16'hcaca;
    LUT4 mux_423_i11_3_lut (.A(quad_count[10]), .B(quad_buffer[10]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i11_3_lut.init = 16'hcaca;
    LUT4 mux_423_i10_3_lut (.A(quad_count[9]), .B(quad_buffer[9]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i10_3_lut.init = 16'hcaca;
    LUT4 mux_423_i9_3_lut (.A(quad_count[8]), .B(quad_buffer[8]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i9_3_lut.init = 16'hcaca;
    LUT4 mux_423_i8_3_lut (.A(quad_count[7]), .B(quad_buffer[7]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i8_3_lut.init = 16'hcaca;
    LUT4 mux_423_i7_3_lut (.A(quad_count[6]), .B(quad_buffer[6]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i7_3_lut.init = 16'hcaca;
    LUT4 mux_423_i6_3_lut (.A(quad_count[5]), .B(quad_buffer[5]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i6_3_lut.init = 16'hcaca;
    LUT4 mux_423_i5_3_lut (.A(quad_count[4]), .B(quad_buffer[4]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i5_3_lut.init = 16'hcaca;
    LUT4 mux_423_i4_3_lut (.A(quad_count[3]), .B(quad_buffer[3]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i4_3_lut.init = 16'hcaca;
    LUT4 mux_423_i3_3_lut (.A(quad_count[2]), .B(quad_buffer[2]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i3_3_lut.init = 16'hcaca;
    LUT4 mux_423_i2_3_lut (.A(quad_count[1]), .B(quad_buffer[1]), .C(n47), 
         .Z(spi_data_out_r_39__N_1318[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_423_i2_3_lut.init = 16'hcaca;
    LUT4 i5497_4_lut (.A(n4129[31]), .B(quad_set[31]), .C(n5715), .D(n1), 
         .Z(n9821)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5497_4_lut.init = 16'hc0ca;
    LUT4 i5495_4_lut (.A(n4129[30]), .B(quad_set[30]), .C(n5715), .D(n1), 
         .Z(n9819)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5495_4_lut.init = 16'hc0ca;
    LUT4 i5493_4_lut (.A(n4129[29]), .B(quad_set[29]), .C(n5715), .D(n1), 
         .Z(n9817)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5493_4_lut.init = 16'hc0ca;
    LUT4 i5491_4_lut (.A(n4129[28]), .B(quad_set[28]), .C(n5715), .D(n1), 
         .Z(n9815)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5491_4_lut.init = 16'hc0ca;
    LUT4 i5489_4_lut (.A(n4129[27]), .B(quad_set[27]), .C(n5715), .D(n1), 
         .Z(n9813)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5489_4_lut.init = 16'hc0ca;
    LUT4 i5487_4_lut (.A(n4129[26]), .B(quad_set[26]), .C(n5715), .D(n1), 
         .Z(n9811)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5487_4_lut.init = 16'hc0ca;
    LUT4 i5485_4_lut (.A(n4129[25]), .B(quad_set[25]), .C(n5715), .D(n1), 
         .Z(n9809)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5485_4_lut.init = 16'hc0ca;
    LUT4 i5483_4_lut (.A(n4129[24]), .B(quad_set[24]), .C(n5715), .D(n1), 
         .Z(n9807)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5483_4_lut.init = 16'hc0ca;
    LUT4 i5481_4_lut (.A(n4129[23]), .B(quad_set[23]), .C(n5715), .D(n1), 
         .Z(n9805)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5481_4_lut.init = 16'hc0ca;
    LUT4 i5479_4_lut (.A(n4129[22]), .B(quad_set[22]), .C(n5715), .D(n1), 
         .Z(n9803)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5479_4_lut.init = 16'hc0ca;
    LUT4 i5477_4_lut (.A(n4129[21]), .B(quad_set[21]), .C(n5715), .D(n1), 
         .Z(n9801)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5477_4_lut.init = 16'hc0ca;
    LUT4 i5475_4_lut (.A(n4129[20]), .B(quad_set[20]), .C(n5715), .D(n1), 
         .Z(n9799)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5475_4_lut.init = 16'hc0ca;
    LUT4 i5473_4_lut (.A(n4129[19]), .B(quad_set[19]), .C(n5715), .D(n1), 
         .Z(n9797)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5473_4_lut.init = 16'hc0ca;
    LUT4 i5471_4_lut (.A(n4129[18]), .B(quad_set[18]), .C(n5715), .D(n1), 
         .Z(n9795)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5471_4_lut.init = 16'hc0ca;
    LUT4 i5469_4_lut (.A(n4129[17]), .B(quad_set[17]), .C(n5715), .D(n1), 
         .Z(n9793)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5469_4_lut.init = 16'hc0ca;
    LUT4 i5467_4_lut (.A(n4129[16]), .B(quad_set[16]), .C(n5715), .D(n1), 
         .Z(n9791)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5467_4_lut.init = 16'hc0ca;
    LUT4 i5465_4_lut (.A(n4129[15]), .B(quad_set[15]), .C(n5715), .D(n1), 
         .Z(n9789)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5465_4_lut.init = 16'hc0ca;
    LUT4 i5463_4_lut (.A(n4129[14]), .B(quad_set[14]), .C(n5715), .D(n1), 
         .Z(n9787)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5463_4_lut.init = 16'hc0ca;
    LUT4 i5461_4_lut (.A(n4129[13]), .B(quad_set[13]), .C(n5715), .D(n1), 
         .Z(n9785)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5461_4_lut.init = 16'hc0ca;
    LUT4 i5459_4_lut (.A(n4129[12]), .B(quad_set[12]), .C(n5715), .D(n1), 
         .Z(n9783)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5459_4_lut.init = 16'hc0ca;
    LUT4 i5457_4_lut (.A(n4129[11]), .B(quad_set[11]), .C(n5715), .D(n1), 
         .Z(n9781)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5457_4_lut.init = 16'hc0ca;
    LUT4 i5455_4_lut (.A(n4129[10]), .B(quad_set[10]), .C(n5715), .D(n1), 
         .Z(n9779)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5455_4_lut.init = 16'hc0ca;
    LUT4 i5453_4_lut (.A(n4129[9]), .B(quad_set[9]), .C(n5715), .D(n1), 
         .Z(n9777)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5453_4_lut.init = 16'hc0ca;
    LUT4 i5451_4_lut (.A(n4129[8]), .B(quad_set[8]), .C(n5715), .D(n1), 
         .Z(n9775)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5451_4_lut.init = 16'hc0ca;
    LUT4 i5449_4_lut (.A(n4129[7]), .B(quad_set[7]), .C(n5715), .D(n1), 
         .Z(n9773)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5449_4_lut.init = 16'hc0ca;
    LUT4 i5447_4_lut (.A(n4129[6]), .B(quad_set[6]), .C(n5715), .D(n1), 
         .Z(n9771)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5447_4_lut.init = 16'hc0ca;
    LUT4 i5445_4_lut (.A(n4129[5]), .B(quad_set[5]), .C(n5715), .D(n1), 
         .Z(n9769)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5445_4_lut.init = 16'hc0ca;
    LUT4 i5443_4_lut (.A(n4129[4]), .B(quad_set[4]), .C(n5715), .D(n1), 
         .Z(n9767)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5443_4_lut.init = 16'hc0ca;
    LUT4 i5441_4_lut (.A(n4129[3]), .B(quad_set[3]), .C(n5715), .D(n1), 
         .Z(n9765)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5441_4_lut.init = 16'hc0ca;
    LUT4 i5439_4_lut (.A(n4129[2]), .B(quad_set[2]), .C(n5715), .D(n1), 
         .Z(n9763)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5439_4_lut.init = 16'hc0ca;
    LUT4 i5437_4_lut (.A(n4129[1]), .B(quad_set[1]), .C(n5715), .D(n1), 
         .Z(n9761)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5437_4_lut.init = 16'hc0ca;
    CCU2D add_1361_33 (.A0(quad_count[30]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[31]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22125), .S0(n4129[30]), .S1(n4129[31]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_33.INIT0 = 16'h5569;
    defparam add_1361_33.INIT1 = 16'h5569;
    defparam add_1361_33.INJECT1_0 = "NO";
    defparam add_1361_33.INJECT1_1 = "NO";
    CCU2D add_1361_31 (.A0(quad_count[28]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[29]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22124), .COUT(n22125), .S0(n4129[28]), .S1(n4129[29]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_31.INIT0 = 16'h5569;
    defparam add_1361_31.INIT1 = 16'h5569;
    defparam add_1361_31.INJECT1_0 = "NO";
    defparam add_1361_31.INJECT1_1 = "NO";
    CCU2D add_1361_29 (.A0(quad_count[26]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[27]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22123), .COUT(n22124), .S0(n4129[26]), .S1(n4129[27]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_29.INIT0 = 16'h5569;
    defparam add_1361_29.INIT1 = 16'h5569;
    defparam add_1361_29.INJECT1_0 = "NO";
    defparam add_1361_29.INJECT1_1 = "NO";
    CCU2D add_1361_27 (.A0(quad_count[24]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[25]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22122), .COUT(n22123), .S0(n4129[24]), .S1(n4129[25]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1361_27.INIT0 = 16'h5569;
    defparam add_1361_27.INIT1 = 16'h5569;
    defparam add_1361_27.INJECT1_0 = "NO";
    defparam add_1361_27.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(quad_homing[0]), .B(quad_homing[1]), .C(quad_set_valid), 
         .D(resetn_c), .Z(n5715)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut.init = 16'h1000;
    LUT4 i24202_2_lut (.A(resetn_c), .B(quad_homing[1]), .Z(clk_enable_519)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i24202_2_lut.init = 16'h7777;
    
endmodule
//
// Verilog Description of module \quad_decoder(DEV_ID=6) 
//

module \quad_decoder(DEV_ID=6)  (GND_net, quad_count, clk, n30185, \quad_a[6] , 
            \quad_b[6] , \spi_data_out_r_39__N_2344[0] , \spi_data_out_r_39__N_2493[0] , 
            quad_buffer, \pin_intrpt[20] , n30004, spi_data_out_r_39__N_2384, 
            spi_data_out_r_39__N_2573, quad_homing, clk_enable_639, \spi_data_r[0] , 
            clk_enable_898, \spi_data_out_r_39__N_2344[31] , \spi_data_out_r_39__N_2493[31] , 
            \spi_data_out_r_39__N_2344[30] , \spi_data_out_r_39__N_2493[30] , 
            \spi_data_out_r_39__N_2344[29] , \spi_data_out_r_39__N_2493[29] , 
            \spi_data_out_r_39__N_2344[28] , \spi_data_out_r_39__N_2493[28] , 
            \spi_data_out_r_39__N_2344[27] , \spi_data_out_r_39__N_2493[27] , 
            \spi_data_out_r_39__N_2344[26] , \spi_data_out_r_39__N_2493[26] , 
            \spi_data_out_r_39__N_2344[25] , \spi_data_out_r_39__N_2493[25] , 
            \spi_data_out_r_39__N_2344[24] , \spi_data_out_r_39__N_2493[24] , 
            \spi_data_out_r_39__N_2344[23] , \spi_data_out_r_39__N_2493[23] , 
            \spi_data_out_r_39__N_2344[22] , \spi_data_out_r_39__N_2493[22] , 
            \spi_data_out_r_39__N_2344[21] , \spi_data_out_r_39__N_2493[21] , 
            \spi_data_out_r_39__N_2344[20] , \spi_data_out_r_39__N_2493[20] , 
            \spi_data_out_r_39__N_2344[19] , \spi_data_out_r_39__N_2493[19] , 
            \spi_data_out_r_39__N_2344[18] , \spi_data_out_r_39__N_2493[18] , 
            \spi_data_out_r_39__N_2344[17] , \spi_data_out_r_39__N_2493[17] , 
            \spi_data_out_r_39__N_2344[16] , \spi_data_out_r_39__N_2493[16] , 
            \spi_data_out_r_39__N_2344[15] , \spi_data_out_r_39__N_2493[15] , 
            \spi_data_out_r_39__N_2344[14] , \spi_data_out_r_39__N_2493[14] , 
            \spi_data_out_r_39__N_2344[13] , \spi_data_out_r_39__N_2493[13] , 
            \spi_data_out_r_39__N_2344[12] , \spi_data_out_r_39__N_2493[12] , 
            \spi_data_out_r_39__N_2344[11] , \spi_data_out_r_39__N_2493[11] , 
            \spi_data_out_r_39__N_2344[10] , \spi_data_out_r_39__N_2493[10] , 
            \spi_data_out_r_39__N_2344[9] , \spi_data_out_r_39__N_2493[9] , 
            \spi_data_out_r_39__N_2344[8] , \spi_data_out_r_39__N_2493[8] , 
            \spi_data_out_r_39__N_2344[7] , \spi_data_out_r_39__N_2493[7] , 
            \spi_data_out_r_39__N_2344[6] , \spi_data_out_r_39__N_2493[6] , 
            \spi_data_out_r_39__N_2344[5] , \spi_data_out_r_39__N_2493[5] , 
            \spi_data_out_r_39__N_2344[4] , \spi_data_out_r_39__N_2493[4] , 
            \spi_data_out_r_39__N_2344[3] , \spi_data_out_r_39__N_2493[3] , 
            \spi_data_out_r_39__N_2344[2] , \spi_data_out_r_39__N_2493[2] , 
            \spi_data_out_r_39__N_2344[1] , \spi_data_out_r_39__N_2493[1] , 
            \spi_data_r[1] , \spi_data_r[2] , \spi_data_r[3] , \spi_data_r[4] , 
            \spi_data_r[5] , \spi_data_r[6] , \spi_data_r[7] , \spi_data_r[8] , 
            \spi_data_r[9] , \spi_data_r[10] , \spi_data_r[11] , \spi_data_r[12] , 
            \spi_data_r[13] , \spi_data_r[14] , \spi_data_r[15] , \spi_data_r[16] , 
            \spi_data_r[17] , \spi_data_r[18] , \spi_data_r[19] , \spi_data_r[20] , 
            \spi_data_r[21] , \spi_data_r[22] , \spi_data_r[23] , \spi_data_r[24] , 
            \spi_data_r[25] , \spi_data_r[26] , \spi_data_r[27] , \spi_data_r[28] , 
            \spi_data_r[29] , \spi_data_r[30] , \spi_data_r[31] , resetn_c, 
            n1) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output [31:0]quad_count;
    input clk;
    input n30185;
    input \quad_a[6] ;
    input \quad_b[6] ;
    output \spi_data_out_r_39__N_2344[0] ;
    input \spi_data_out_r_39__N_2493[0] ;
    output [31:0]quad_buffer;
    input \pin_intrpt[20] ;
    input n30004;
    output spi_data_out_r_39__N_2384;
    input spi_data_out_r_39__N_2573;
    output [1:0]quad_homing;
    input clk_enable_639;
    input \spi_data_r[0] ;
    input clk_enable_898;
    output \spi_data_out_r_39__N_2344[31] ;
    input \spi_data_out_r_39__N_2493[31] ;
    output \spi_data_out_r_39__N_2344[30] ;
    input \spi_data_out_r_39__N_2493[30] ;
    output \spi_data_out_r_39__N_2344[29] ;
    input \spi_data_out_r_39__N_2493[29] ;
    output \spi_data_out_r_39__N_2344[28] ;
    input \spi_data_out_r_39__N_2493[28] ;
    output \spi_data_out_r_39__N_2344[27] ;
    input \spi_data_out_r_39__N_2493[27] ;
    output \spi_data_out_r_39__N_2344[26] ;
    input \spi_data_out_r_39__N_2493[26] ;
    output \spi_data_out_r_39__N_2344[25] ;
    input \spi_data_out_r_39__N_2493[25] ;
    output \spi_data_out_r_39__N_2344[24] ;
    input \spi_data_out_r_39__N_2493[24] ;
    output \spi_data_out_r_39__N_2344[23] ;
    input \spi_data_out_r_39__N_2493[23] ;
    output \spi_data_out_r_39__N_2344[22] ;
    input \spi_data_out_r_39__N_2493[22] ;
    output \spi_data_out_r_39__N_2344[21] ;
    input \spi_data_out_r_39__N_2493[21] ;
    output \spi_data_out_r_39__N_2344[20] ;
    input \spi_data_out_r_39__N_2493[20] ;
    output \spi_data_out_r_39__N_2344[19] ;
    input \spi_data_out_r_39__N_2493[19] ;
    output \spi_data_out_r_39__N_2344[18] ;
    input \spi_data_out_r_39__N_2493[18] ;
    output \spi_data_out_r_39__N_2344[17] ;
    input \spi_data_out_r_39__N_2493[17] ;
    output \spi_data_out_r_39__N_2344[16] ;
    input \spi_data_out_r_39__N_2493[16] ;
    output \spi_data_out_r_39__N_2344[15] ;
    input \spi_data_out_r_39__N_2493[15] ;
    output \spi_data_out_r_39__N_2344[14] ;
    input \spi_data_out_r_39__N_2493[14] ;
    output \spi_data_out_r_39__N_2344[13] ;
    input \spi_data_out_r_39__N_2493[13] ;
    output \spi_data_out_r_39__N_2344[12] ;
    input \spi_data_out_r_39__N_2493[12] ;
    output \spi_data_out_r_39__N_2344[11] ;
    input \spi_data_out_r_39__N_2493[11] ;
    output \spi_data_out_r_39__N_2344[10] ;
    input \spi_data_out_r_39__N_2493[10] ;
    output \spi_data_out_r_39__N_2344[9] ;
    input \spi_data_out_r_39__N_2493[9] ;
    output \spi_data_out_r_39__N_2344[8] ;
    input \spi_data_out_r_39__N_2493[8] ;
    output \spi_data_out_r_39__N_2344[7] ;
    input \spi_data_out_r_39__N_2493[7] ;
    output \spi_data_out_r_39__N_2344[6] ;
    input \spi_data_out_r_39__N_2493[6] ;
    output \spi_data_out_r_39__N_2344[5] ;
    input \spi_data_out_r_39__N_2493[5] ;
    output \spi_data_out_r_39__N_2344[4] ;
    input \spi_data_out_r_39__N_2493[4] ;
    output \spi_data_out_r_39__N_2344[3] ;
    input \spi_data_out_r_39__N_2493[3] ;
    output \spi_data_out_r_39__N_2344[2] ;
    input \spi_data_out_r_39__N_2493[2] ;
    output \spi_data_out_r_39__N_2344[1] ;
    input \spi_data_out_r_39__N_2493[1] ;
    input \spi_data_r[1] ;
    input \spi_data_r[2] ;
    input \spi_data_r[3] ;
    input \spi_data_r[4] ;
    input \spi_data_r[5] ;
    input \spi_data_r[6] ;
    input \spi_data_r[7] ;
    input \spi_data_r[8] ;
    input \spi_data_r[9] ;
    input \spi_data_r[10] ;
    input \spi_data_r[11] ;
    input \spi_data_r[12] ;
    input \spi_data_r[13] ;
    input \spi_data_r[14] ;
    input \spi_data_r[15] ;
    input \spi_data_r[16] ;
    input \spi_data_r[17] ;
    input \spi_data_r[18] ;
    input \spi_data_r[19] ;
    input \spi_data_r[20] ;
    input \spi_data_r[21] ;
    input \spi_data_r[22] ;
    input \spi_data_r[23] ;
    input \spi_data_r[24] ;
    input \spi_data_r[25] ;
    input \spi_data_r[26] ;
    input \spi_data_r[27] ;
    input \spi_data_r[28] ;
    input \spi_data_r[29] ;
    input \spi_data_r[30] ;
    input \spi_data_r[31] ;
    input resetn_c;
    input n1;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire \pin_intrpt[20]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[20] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    wire [2:0]quad_a_delayed;   // c:/s_links/sources/quad_decoder.v(34[20:34])
    wire [2:0]quad_b_delayed;   // c:/s_links/sources/quad_decoder.v(35[19:33])
    
    wire n21997, clk_enable_353, n7967, quad_set_valid;
    wire [31:0]quad_set;   // c:/s_links/sources/quad_decoder.v(39[31:39])
    
    wire n8716, n8718, n8720, n8722, n8724, n8726, n8728, n8730, 
        n8732, n8734, n8736, n8738, n8740, n8742, n8744, n8772, 
        n8774, n8776, n8778, n8780, n8782, n8784, n8786, n8788, 
        n8790, n8792, n8794, n8796, n8798, n8800, n8802, n6, 
        count_dir, n22012;
    wire [31:0]n4096;
    
    wire n22011, n22010, n22009, n22008, n22007, n5695, n22006, 
        n22005, n22004, n22003, n22002, n22001, n22000, n21999, 
        n21998;
    
    CCU2D add_1377_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quad_a_delayed[2]), .B1(quad_b_delayed[1]), .C1(quad_b_delayed[2]), 
          .D1(quad_a_delayed[1]), .COUT(n21997));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_1.INIT0 = 16'hF000;
    defparam add_1377_1.INIT1 = 16'h0990;
    defparam add_1377_1.INJECT1_0 = "NO";
    defparam add_1377_1.INJECT1_1 = "NO";
    FD1P3AX quad_count_i0_i0 (.D(n7967), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i0.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i0 (.D(\quad_a[6] ), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i0.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i0 (.D(\quad_b[6] ), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_2493[0] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX quad_buffer_i0 (.D(quad_count[0]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i0.GSR = "DISABLED";
    FD1S3IX quad_set_valid_388 (.D(n30004), .CK(clk), .CD(n30185), .Q(quad_set_valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set_valid_388.GSR = "DISABLED";
    FD1S3IX i39_391 (.D(spi_data_out_r_39__N_2573), .CK(clk), .CD(n30185), 
            .Q(spi_data_out_r_39__N_2384)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam i39_391.GSR = "DISABLED";
    FD1P3IX quad_homing__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_639), .CD(n30185), 
            .CK(clk), .Q(quad_homing[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(62[8] 69[4])
    defparam quad_homing__i0.GSR = "DISABLED";
    FD1P3IX quad_set__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i0.GSR = "DISABLED";
    FD1S3AX quad_buffer_i31 (.D(quad_count[31]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i31.GSR = "DISABLED";
    FD1S3AX quad_buffer_i30 (.D(quad_count[30]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i30.GSR = "DISABLED";
    FD1S3AX quad_buffer_i29 (.D(quad_count[29]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i29.GSR = "DISABLED";
    FD1S3AX quad_buffer_i28 (.D(quad_count[28]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i28.GSR = "DISABLED";
    FD1S3AX quad_buffer_i27 (.D(quad_count[27]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i27.GSR = "DISABLED";
    FD1S3AX quad_buffer_i26 (.D(quad_count[26]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i26.GSR = "DISABLED";
    FD1S3AX quad_buffer_i25 (.D(quad_count[25]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i25.GSR = "DISABLED";
    FD1S3AX quad_buffer_i24 (.D(quad_count[24]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i24.GSR = "DISABLED";
    FD1S3AX quad_buffer_i23 (.D(quad_count[23]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i23.GSR = "DISABLED";
    FD1S3AX quad_buffer_i22 (.D(quad_count[22]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i22.GSR = "DISABLED";
    FD1S3AX quad_buffer_i21 (.D(quad_count[21]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i21.GSR = "DISABLED";
    FD1S3AX quad_buffer_i20 (.D(quad_count[20]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i20.GSR = "DISABLED";
    FD1S3AX quad_buffer_i19 (.D(quad_count[19]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i19.GSR = "DISABLED";
    FD1S3AX quad_buffer_i18 (.D(quad_count[18]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i18.GSR = "DISABLED";
    FD1S3AX quad_buffer_i17 (.D(quad_count[17]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i17.GSR = "DISABLED";
    FD1S3AX quad_buffer_i16 (.D(quad_count[16]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i16.GSR = "DISABLED";
    FD1S3AX quad_buffer_i15 (.D(quad_count[15]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i15.GSR = "DISABLED";
    FD1S3AX quad_buffer_i14 (.D(quad_count[14]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i14.GSR = "DISABLED";
    FD1S3AX quad_buffer_i13 (.D(quad_count[13]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i13.GSR = "DISABLED";
    FD1S3AX quad_buffer_i12 (.D(quad_count[12]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i12.GSR = "DISABLED";
    FD1S3AX quad_buffer_i11 (.D(quad_count[11]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i11.GSR = "DISABLED";
    FD1S3AX quad_buffer_i10 (.D(quad_count[10]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i10.GSR = "DISABLED";
    FD1S3AX quad_buffer_i9 (.D(quad_count[9]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i9.GSR = "DISABLED";
    FD1S3AX quad_buffer_i8 (.D(quad_count[8]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i8.GSR = "DISABLED";
    FD1S3AX quad_buffer_i7 (.D(quad_count[7]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i7.GSR = "DISABLED";
    FD1S3AX quad_buffer_i6 (.D(quad_count[6]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i6.GSR = "DISABLED";
    FD1S3AX quad_buffer_i5 (.D(quad_count[5]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i5.GSR = "DISABLED";
    FD1S3AX quad_buffer_i4 (.D(quad_count[4]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i4.GSR = "DISABLED";
    FD1S3AX quad_buffer_i3 (.D(quad_count[3]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i3.GSR = "DISABLED";
    FD1S3AX quad_buffer_i2 (.D(quad_count[2]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i2.GSR = "DISABLED";
    FD1S3AX quad_buffer_i1 (.D(quad_count[1]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_2493[31] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i31 (.D(\spi_data_out_r_39__N_2493[30] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i30 (.D(\spi_data_out_r_39__N_2493[29] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i29 (.D(\spi_data_out_r_39__N_2493[28] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i28 (.D(\spi_data_out_r_39__N_2493[27] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i27 (.D(\spi_data_out_r_39__N_2493[26] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i26 (.D(\spi_data_out_r_39__N_2493[25] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i25 (.D(\spi_data_out_r_39__N_2493[24] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i24 (.D(\spi_data_out_r_39__N_2493[23] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i23 (.D(\spi_data_out_r_39__N_2493[22] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i22 (.D(\spi_data_out_r_39__N_2493[21] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i21 (.D(\spi_data_out_r_39__N_2493[20] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i20 (.D(\spi_data_out_r_39__N_2493[19] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i19 (.D(\spi_data_out_r_39__N_2493[18] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i18 (.D(\spi_data_out_r_39__N_2493[17] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i17 (.D(\spi_data_out_r_39__N_2493[16] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i16 (.D(\spi_data_out_r_39__N_2493[15] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_2493[14] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_2493[13] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_2493[12] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_2493[11] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_2493[10] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_2493[9] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_2493[8] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_2493[7] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_2493[6] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_2493[5] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_2493[4] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_2493[3] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_2493[2] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_2493[1] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2344[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i2 (.D(quad_b_delayed[1]), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i2.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i1 (.D(quad_b_delayed[0]), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i1.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i2 (.D(quad_a_delayed[1]), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i2.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i1 (.D(quad_a_delayed[0]), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i1.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i31 (.D(n8716), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i31.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i30 (.D(n8718), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i30.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i29 (.D(n8720), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i29.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i28 (.D(n8722), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i28.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i27 (.D(n8724), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i27.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i26 (.D(n8726), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i26.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i25 (.D(n8728), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i25.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i24 (.D(n8730), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i24.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i23 (.D(n8732), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i23.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i22 (.D(n8734), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i22.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i21 (.D(n8736), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i21.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i20 (.D(n8738), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i20.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i19 (.D(n8740), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i19.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i18 (.D(n8742), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i18.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i17 (.D(n8744), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i17.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i16 (.D(n8772), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i16.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i15 (.D(n8774), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i15.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i14 (.D(n8776), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i14.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i13 (.D(n8778), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i13.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i12 (.D(n8780), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i12.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i11 (.D(n8782), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i11.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i10 (.D(n8784), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i10.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i9 (.D(n8786), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i9.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i8 (.D(n8788), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i8.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i7 (.D(n8790), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i7.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i6 (.D(n8792), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i6.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i5 (.D(n8794), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i5.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i4 (.D(n8796), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i4.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i3 (.D(n8798), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i3.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i2 (.D(n8800), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i1 (.D(n8802), .SP(clk_enable_353), .CK(clk), 
            .Q(quad_count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i1.GSR = "DISABLED";
    FD1P3IX quad_homing__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_639), .CD(n30185), 
            .CK(clk), .Q(quad_homing[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(62[8] 69[4])
    defparam quad_homing__i1.GSR = "DISABLED";
    LUT4 i2_2_lut (.A(quad_b_delayed[1]), .B(quad_a_delayed[2]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(96[19:96])
    defparam i2_2_lut.init = 16'h6666;
    LUT4 i1_2_lut (.A(quad_a_delayed[1]), .B(quad_b_delayed[2]), .Z(count_dir)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(96[19:96])
    defparam i1_2_lut.init = 16'h6666;
    FD1P3IX quad_set__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i1.GSR = "DISABLED";
    FD1P3IX quad_set__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i2.GSR = "DISABLED";
    FD1P3IX quad_set__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i3.GSR = "DISABLED";
    FD1P3IX quad_set__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i4.GSR = "DISABLED";
    FD1P3IX quad_set__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i5.GSR = "DISABLED";
    FD1P3IX quad_set__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i6.GSR = "DISABLED";
    FD1P3IX quad_set__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i7.GSR = "DISABLED";
    FD1P3IX quad_set__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i8.GSR = "DISABLED";
    FD1P3IX quad_set__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i9.GSR = "DISABLED";
    FD1P3IX quad_set__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i10.GSR = "DISABLED";
    FD1P3IX quad_set__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i11.GSR = "DISABLED";
    FD1P3IX quad_set__i12 (.D(\spi_data_r[12] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i12.GSR = "DISABLED";
    FD1P3IX quad_set__i13 (.D(\spi_data_r[13] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i13.GSR = "DISABLED";
    FD1P3IX quad_set__i14 (.D(\spi_data_r[14] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i14.GSR = "DISABLED";
    FD1P3IX quad_set__i15 (.D(\spi_data_r[15] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i15.GSR = "DISABLED";
    FD1P3IX quad_set__i16 (.D(\spi_data_r[16] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i16.GSR = "DISABLED";
    FD1P3IX quad_set__i17 (.D(\spi_data_r[17] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i17.GSR = "DISABLED";
    FD1P3IX quad_set__i18 (.D(\spi_data_r[18] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i18.GSR = "DISABLED";
    FD1P3IX quad_set__i19 (.D(\spi_data_r[19] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i19.GSR = "DISABLED";
    FD1P3IX quad_set__i20 (.D(\spi_data_r[20] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i20.GSR = "DISABLED";
    FD1P3IX quad_set__i21 (.D(\spi_data_r[21] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i21.GSR = "DISABLED";
    FD1P3IX quad_set__i22 (.D(\spi_data_r[22] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i22.GSR = "DISABLED";
    FD1P3IX quad_set__i23 (.D(\spi_data_r[23] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i23.GSR = "DISABLED";
    FD1P3IX quad_set__i24 (.D(\spi_data_r[24] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i24.GSR = "DISABLED";
    FD1P3IX quad_set__i25 (.D(\spi_data_r[25] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i25.GSR = "DISABLED";
    FD1P3IX quad_set__i26 (.D(\spi_data_r[26] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i26.GSR = "DISABLED";
    FD1P3IX quad_set__i27 (.D(\spi_data_r[27] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i27.GSR = "DISABLED";
    FD1P3IX quad_set__i28 (.D(\spi_data_r[28] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i28.GSR = "DISABLED";
    FD1P3IX quad_set__i29 (.D(\spi_data_r[29] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i29.GSR = "DISABLED";
    FD1P3IX quad_set__i30 (.D(\spi_data_r[30] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i30.GSR = "DISABLED";
    FD1P3IX quad_set__i31 (.D(\spi_data_r[31] ), .SP(clk_enable_898), .CD(n30185), 
            .CK(clk), .Q(quad_set[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i31.GSR = "DISABLED";
    CCU2D add_1377_33 (.A0(quad_count[30]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[31]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22012), .S0(n4096[30]), .S1(n4096[31]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_33.INIT0 = 16'h5569;
    defparam add_1377_33.INIT1 = 16'h5569;
    defparam add_1377_33.INJECT1_0 = "NO";
    defparam add_1377_33.INJECT1_1 = "NO";
    CCU2D add_1377_31 (.A0(quad_count[28]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[29]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22011), .COUT(n22012), .S0(n4096[28]), .S1(n4096[29]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_31.INIT0 = 16'h5569;
    defparam add_1377_31.INIT1 = 16'h5569;
    defparam add_1377_31.INJECT1_0 = "NO";
    defparam add_1377_31.INJECT1_1 = "NO";
    CCU2D add_1377_29 (.A0(quad_count[26]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[27]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22010), .COUT(n22011), .S0(n4096[26]), .S1(n4096[27]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_29.INIT0 = 16'h5569;
    defparam add_1377_29.INIT1 = 16'h5569;
    defparam add_1377_29.INJECT1_0 = "NO";
    defparam add_1377_29.INJECT1_1 = "NO";
    CCU2D add_1377_27 (.A0(quad_count[24]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[25]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22009), .COUT(n22010), .S0(n4096[24]), .S1(n4096[25]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_27.INIT0 = 16'h5569;
    defparam add_1377_27.INIT1 = 16'h5569;
    defparam add_1377_27.INJECT1_0 = "NO";
    defparam add_1377_27.INJECT1_1 = "NO";
    LUT4 i24181_2_lut (.A(resetn_c), .B(quad_homing[1]), .Z(clk_enable_353)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i24181_2_lut.init = 16'h7777;
    CCU2D add_1377_25 (.A0(quad_count[22]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[23]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22008), .COUT(n22009), .S0(n4096[22]), .S1(n4096[23]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_25.INIT0 = 16'h5569;
    defparam add_1377_25.INIT1 = 16'h5569;
    defparam add_1377_25.INJECT1_0 = "NO";
    defparam add_1377_25.INJECT1_1 = "NO";
    CCU2D add_1377_23 (.A0(quad_count[20]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[21]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22007), .COUT(n22008), .S0(n4096[20]), .S1(n4096[21]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_23.INIT0 = 16'h5569;
    defparam add_1377_23.INIT1 = 16'h5569;
    defparam add_1377_23.INJECT1_0 = "NO";
    defparam add_1377_23.INJECT1_1 = "NO";
    LUT4 i3645_4_lut (.A(n4096[0]), .B(quad_set[0]), .C(n5695), .D(n1), 
         .Z(n7967)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i3645_4_lut.init = 16'hc0ca;
    LUT4 i1_4_lut (.A(quad_homing[0]), .B(quad_homing[1]), .C(quad_set_valid), 
         .D(resetn_c), .Z(n5695)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut.init = 16'h1000;
    CCU2D add_1377_21 (.A0(quad_count[18]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[19]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22006), .COUT(n22007), .S0(n4096[18]), .S1(n4096[19]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_21.INIT0 = 16'h5569;
    defparam add_1377_21.INIT1 = 16'h5569;
    defparam add_1377_21.INJECT1_0 = "NO";
    defparam add_1377_21.INJECT1_1 = "NO";
    CCU2D add_1377_19 (.A0(quad_count[16]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[17]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22005), .COUT(n22006), .S0(n4096[16]), .S1(n4096[17]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_19.INIT0 = 16'h5569;
    defparam add_1377_19.INIT1 = 16'h5569;
    defparam add_1377_19.INJECT1_0 = "NO";
    defparam add_1377_19.INJECT1_1 = "NO";
    CCU2D add_1377_17 (.A0(quad_count[14]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[15]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22004), .COUT(n22005), .S0(n4096[14]), .S1(n4096[15]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_17.INIT0 = 16'h5569;
    defparam add_1377_17.INIT1 = 16'h5569;
    defparam add_1377_17.INJECT1_0 = "NO";
    defparam add_1377_17.INJECT1_1 = "NO";
    CCU2D add_1377_15 (.A0(quad_count[12]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[13]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22003), .COUT(n22004), .S0(n4096[12]), .S1(n4096[13]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_15.INIT0 = 16'h5569;
    defparam add_1377_15.INIT1 = 16'h5569;
    defparam add_1377_15.INJECT1_0 = "NO";
    defparam add_1377_15.INJECT1_1 = "NO";
    CCU2D add_1377_13 (.A0(quad_count[10]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[11]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22002), .COUT(n22003), .S0(n4096[10]), .S1(n4096[11]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_13.INIT0 = 16'h5569;
    defparam add_1377_13.INIT1 = 16'h5569;
    defparam add_1377_13.INJECT1_0 = "NO";
    defparam add_1377_13.INJECT1_1 = "NO";
    CCU2D add_1377_11 (.A0(quad_count[8]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[9]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22001), .COUT(n22002), .S0(n4096[8]), .S1(n4096[9]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_11.INIT0 = 16'h5569;
    defparam add_1377_11.INIT1 = 16'h5569;
    defparam add_1377_11.INJECT1_0 = "NO";
    defparam add_1377_11.INJECT1_1 = "NO";
    LUT4 i4392_4_lut (.A(n4096[31]), .B(quad_set[31]), .C(n5695), .D(n1), 
         .Z(n8716)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4392_4_lut.init = 16'hc0ca;
    CCU2D add_1377_9 (.A0(quad_count[6]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[7]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22000), .COUT(n22001), .S0(n4096[6]), .S1(n4096[7]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_9.INIT0 = 16'h5569;
    defparam add_1377_9.INIT1 = 16'h5569;
    defparam add_1377_9.INJECT1_0 = "NO";
    defparam add_1377_9.INJECT1_1 = "NO";
    LUT4 i4394_4_lut (.A(n4096[30]), .B(quad_set[30]), .C(n5695), .D(n1), 
         .Z(n8718)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4394_4_lut.init = 16'hc0ca;
    CCU2D add_1377_7 (.A0(quad_count[4]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[5]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21999), .COUT(n22000), .S0(n4096[4]), .S1(n4096[5]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_7.INIT0 = 16'h5569;
    defparam add_1377_7.INIT1 = 16'h5569;
    defparam add_1377_7.INJECT1_0 = "NO";
    defparam add_1377_7.INJECT1_1 = "NO";
    LUT4 i4396_4_lut (.A(n4096[29]), .B(quad_set[29]), .C(n5695), .D(n1), 
         .Z(n8720)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4396_4_lut.init = 16'hc0ca;
    LUT4 i4398_4_lut (.A(n4096[28]), .B(quad_set[28]), .C(n5695), .D(n1), 
         .Z(n8722)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4398_4_lut.init = 16'hc0ca;
    LUT4 i4400_4_lut (.A(n4096[27]), .B(quad_set[27]), .C(n5695), .D(n1), 
         .Z(n8724)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4400_4_lut.init = 16'hc0ca;
    LUT4 i4402_4_lut (.A(n4096[26]), .B(quad_set[26]), .C(n5695), .D(n1), 
         .Z(n8726)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4402_4_lut.init = 16'hc0ca;
    LUT4 i4404_4_lut (.A(n4096[25]), .B(quad_set[25]), .C(n5695), .D(n1), 
         .Z(n8728)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4404_4_lut.init = 16'hc0ca;
    LUT4 i4406_4_lut (.A(n4096[24]), .B(quad_set[24]), .C(n5695), .D(n1), 
         .Z(n8730)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4406_4_lut.init = 16'hc0ca;
    LUT4 i4408_4_lut (.A(n4096[23]), .B(quad_set[23]), .C(n5695), .D(n1), 
         .Z(n8732)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4408_4_lut.init = 16'hc0ca;
    LUT4 i4410_4_lut (.A(n4096[22]), .B(quad_set[22]), .C(n5695), .D(n1), 
         .Z(n8734)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4410_4_lut.init = 16'hc0ca;
    LUT4 i4412_4_lut (.A(n4096[21]), .B(quad_set[21]), .C(n5695), .D(n1), 
         .Z(n8736)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4412_4_lut.init = 16'hc0ca;
    LUT4 i4414_4_lut (.A(n4096[20]), .B(quad_set[20]), .C(n5695), .D(n1), 
         .Z(n8738)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4414_4_lut.init = 16'hc0ca;
    LUT4 i4416_4_lut (.A(n4096[19]), .B(quad_set[19]), .C(n5695), .D(n1), 
         .Z(n8740)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4416_4_lut.init = 16'hc0ca;
    LUT4 i4418_4_lut (.A(n4096[18]), .B(quad_set[18]), .C(n5695), .D(n1), 
         .Z(n8742)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4418_4_lut.init = 16'hc0ca;
    LUT4 i4420_4_lut (.A(n4096[17]), .B(quad_set[17]), .C(n5695), .D(n1), 
         .Z(n8744)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4420_4_lut.init = 16'hc0ca;
    LUT4 i4448_4_lut (.A(n4096[16]), .B(quad_set[16]), .C(n5695), .D(n1), 
         .Z(n8772)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4448_4_lut.init = 16'hc0ca;
    LUT4 i4450_4_lut (.A(n4096[15]), .B(quad_set[15]), .C(n5695), .D(n1), 
         .Z(n8774)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4450_4_lut.init = 16'hc0ca;
    LUT4 i4452_4_lut (.A(n4096[14]), .B(quad_set[14]), .C(n5695), .D(n1), 
         .Z(n8776)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4452_4_lut.init = 16'hc0ca;
    LUT4 i4454_4_lut (.A(n4096[13]), .B(quad_set[13]), .C(n5695), .D(n1), 
         .Z(n8778)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4454_4_lut.init = 16'hc0ca;
    LUT4 i4456_4_lut (.A(n4096[12]), .B(quad_set[12]), .C(n5695), .D(n1), 
         .Z(n8780)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4456_4_lut.init = 16'hc0ca;
    LUT4 i4458_4_lut (.A(n4096[11]), .B(quad_set[11]), .C(n5695), .D(n1), 
         .Z(n8782)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4458_4_lut.init = 16'hc0ca;
    LUT4 i4460_4_lut (.A(n4096[10]), .B(quad_set[10]), .C(n5695), .D(n1), 
         .Z(n8784)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4460_4_lut.init = 16'hc0ca;
    LUT4 i4462_4_lut (.A(n4096[9]), .B(quad_set[9]), .C(n5695), .D(n1), 
         .Z(n8786)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4462_4_lut.init = 16'hc0ca;
    LUT4 i4464_4_lut (.A(n4096[8]), .B(quad_set[8]), .C(n5695), .D(n1), 
         .Z(n8788)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4464_4_lut.init = 16'hc0ca;
    LUT4 i4466_4_lut (.A(n4096[7]), .B(quad_set[7]), .C(n5695), .D(n1), 
         .Z(n8790)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4466_4_lut.init = 16'hc0ca;
    LUT4 i4468_4_lut (.A(n4096[6]), .B(quad_set[6]), .C(n5695), .D(n1), 
         .Z(n8792)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4468_4_lut.init = 16'hc0ca;
    LUT4 i4470_4_lut (.A(n4096[5]), .B(quad_set[5]), .C(n5695), .D(n1), 
         .Z(n8794)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4470_4_lut.init = 16'hc0ca;
    LUT4 i4472_4_lut (.A(n4096[4]), .B(quad_set[4]), .C(n5695), .D(n1), 
         .Z(n8796)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4472_4_lut.init = 16'hc0ca;
    LUT4 i4474_4_lut (.A(n4096[3]), .B(quad_set[3]), .C(n5695), .D(n1), 
         .Z(n8798)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4474_4_lut.init = 16'hc0ca;
    LUT4 i4476_4_lut (.A(n4096[2]), .B(quad_set[2]), .C(n5695), .D(n1), 
         .Z(n8800)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4476_4_lut.init = 16'hc0ca;
    LUT4 i4478_4_lut (.A(n4096[1]), .B(quad_set[1]), .C(n5695), .D(n1), 
         .Z(n8802)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4478_4_lut.init = 16'hc0ca;
    CCU2D add_1377_5 (.A0(quad_count[2]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[3]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21998), .COUT(n21999), .S0(n4096[2]), .S1(n4096[3]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_5.INIT0 = 16'h5569;
    defparam add_1377_5.INIT1 = 16'h5569;
    defparam add_1377_5.INJECT1_0 = "NO";
    defparam add_1377_5.INJECT1_1 = "NO";
    CCU2D add_1377_3 (.A0(quad_count[0]), .B0(count_dir), .C0(n6), .D0(count_dir), 
          .A1(quad_count[1]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21997), .COUT(n21998), .S0(n4096[0]), .S1(n4096[1]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1377_3.INIT0 = 16'h5665;
    defparam add_1377_3.INIT1 = 16'h5569;
    defparam add_1377_3.INJECT1_0 = "NO";
    defparam add_1377_3.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \peizo_elliptec(DEV_ID=7,UART_ADDRESS_WIDTH=4) 
//

module \peizo_elliptec(DEV_ID=7,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_32, 
            n30185, \spi_data_r[0] , n28, n29594, uart_slot_en, n30118, 
            n6, n29944, n29943, \spi_cmd_r[0] , spi_addr_r, n30138, 
            \spi_cmd_r[2] , n30023, n26107, n30090, n29481, n25941, 
            n25923, n30062, n30087, pin_io_out_55, n28358, pin_io_out_40, 
            n30122, n24700, n23248, n10696, tx_N_6586, n25358, n30083, 
            mode_adj_656, C_8_c, n30064, n30155, n26091, n30214, 
            n28402, n30094, n28486, n18440, n26113, n26119, n30095, 
            pin_io_out_25, mode_adj_657, n30043, n4, pin_io_out_6, 
            mode_adj_658, mode_adj_659, pin_io_out_5, n30120, n23409, 
            n26089, n25739, n25741) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_32;
    input n30185;
    input \spi_data_r[0] ;
    input n28;
    input n29594;
    input [3:0]uart_slot_en;
    input n30118;
    output n6;
    input n29944;
    input n29943;
    input \spi_cmd_r[0] ;
    input [7:0]spi_addr_r;
    output n30138;
    input \spi_cmd_r[2] ;
    output n30023;
    output n26107;
    output n30090;
    input n29481;
    input n25941;
    output n25923;
    output n30062;
    input n30087;
    input pin_io_out_55;
    output n28358;
    input pin_io_out_40;
    output n30122;
    input n24700;
    output n23248;
    input n10696;
    input tx_N_6586;
    output n25358;
    input n30083;
    input mode_adj_656;
    input C_8_c;
    input n30064;
    input n30155;
    output n26091;
    output n30214;
    output n28402;
    output n30094;
    output n28486;
    input n18440;
    input n26113;
    output n26119;
    input n30095;
    input pin_io_out_25;
    input mode_adj_657;
    input n30043;
    input n4;
    input pin_io_out_6;
    input mode_adj_658;
    input mode_adj_659;
    input pin_io_out_5;
    output n30120;
    output n23409;
    output n26089;
    input n25739;
    output n25741;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    
    wire n29986, n29945, n29984, n29946, n24734, n29485, n29486, 
        n29482, n29483, n29940, n29592, n31066, n29487, n4_c, 
        n29591, n26111, n29590, n52;
    
    FD1P3IX mode_26 (.D(\spi_data_r[0] ), .SP(clk_enable_32), .CD(n30185), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=591, LSE_RLINE=611 */ ;   // c:/s_links/sources/slot_cards/peizo_elliptec.v(36[8] 44[4])
    defparam mode_26.GSR = "DISABLED";
    LUT4 n28_bdd_4_lut_24459 (.A(n28), .B(n29594), .C(uart_slot_en[1]), 
         .D(uart_slot_en[3]), .Z(n29986)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n28_bdd_4_lut_24459.init = 16'hca00;
    LUT4 i1_2_lut_4_lut (.A(uart_slot_en[1]), .B(uart_slot_en[2]), .C(n30118), 
         .D(uart_slot_en[0]), .Z(n6)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h4000;
    L6MUX21 i24385 (.D0(n29945), .D1(n29984), .SD(uart_slot_en[2]), .Z(n29946));
    PFUMX i24383 (.BLUT(n29944), .ALUT(n29943), .C0(uart_slot_en[1]), 
          .Z(n29945));
    LUT4 i1_2_lut_rep_738 (.A(\spi_cmd_r[0] ), .B(spi_addr_r[1]), .Z(n30138)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_738.init = 16'h8888;
    LUT4 i1_2_lut_rep_623_3_lut_4_lut (.A(\spi_cmd_r[0] ), .B(spi_addr_r[1]), 
         .C(spi_addr_r[3]), .D(\spi_cmd_r[2] ), .Z(n30023)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_rep_623_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut (.A(spi_addr_r[3]), .B(spi_addr_r[4]), .Z(n26107)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_rep_690_3_lut (.A(\spi_cmd_r[0] ), .B(spi_addr_r[1]), 
         .C(\spi_cmd_r[2] ), .Z(n30090)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_690_3_lut.init = 16'h8080;
    PFUMX i24238 (.BLUT(n24734), .ALUT(n29485), .C0(uart_slot_en[2]), 
          .Z(n29486));
    PFUMX i24236 (.BLUT(n29482), .ALUT(n29481), .C0(uart_slot_en[3]), 
          .Z(n29483));
    LUT4 i1_2_lut_3_lut_4_lut (.A(\spi_cmd_r[0] ), .B(spi_addr_r[1]), .C(n25941), 
         .D(\spi_cmd_r[2] ), .Z(n25923)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_662_3_lut (.A(\spi_cmd_r[0] ), .B(spi_addr_r[1]), 
         .C(\spi_cmd_r[2] ), .Z(n30062)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_662_3_lut.init = 16'h0808;
    LUT4 RESET_N_5832_bdd_4_lut (.A(n30087), .B(pin_io_out_55), .C(n29940), 
         .D(uart_slot_en[1]), .Z(n29984)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;
    defparam RESET_N_5832_bdd_4_lut.init = 16'hf088;
    LUT4 i23656_2_lut (.A(spi_addr_r[2]), .B(spi_addr_r[4]), .Z(n28358)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23656_2_lut.init = 16'heeee;
    LUT4 n29592_bdd_4_lut (.A(n29592), .B(uart_slot_en[3]), .C(n29986), 
         .D(uart_slot_en[2]), .Z(n31066)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C))) */ ;
    defparam n29592_bdd_4_lut.init = 16'h22f0;
    LUT4 n24734_bdd_3_lut_4_lut (.A(pin_io_out_40), .B(n30122), .C(uart_slot_en[0]), 
         .D(n24700), .Z(n29485)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam n24734_bdd_3_lut_4_lut.init = 16'hf808;
    LUT4 i1_4_lut (.A(uart_slot_en[3]), .B(n29487), .C(n29946), .D(uart_slot_en[0]), 
         .Z(n23248)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'hccec;
    LUT4 i24042_4_lut (.A(n10696), .B(n31066), .C(tx_N_6586), .D(n4_c), 
         .Z(n25358)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+!(C)))) */ ;
    defparam i24042_4_lut.init = 16'h1030;
    LUT4 n29486_bdd_3_lut_4_lut (.A(n29486), .B(n29483), .C(uart_slot_en[0]), 
         .D(uart_slot_en[1]), .Z(n29487)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (C (D)))) */ ;
    defparam n29486_bdd_3_lut_4_lut.init = 16'hc0aa;
    LUT4 i1_4_lut_adj_890 (.A(n30087), .B(uart_slot_en[1]), .C(n30083), 
         .D(uart_slot_en[0]), .Z(n4_c)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_890.init = 16'h3022;
    LUT4 n23552_bdd_2_lut_24364 (.A(mode_adj_656), .B(uart_slot_en[0]), 
         .Z(n29591)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n23552_bdd_2_lut_24364.init = 16'h2222;
    LUT4 RESET_N_5832_bdd_2_lut_24379 (.A(mode), .B(C_8_c), .Z(n29940)) /* synthesis lut_function=(A (B)) */ ;
    defparam RESET_N_5832_bdd_2_lut_24379.init = 16'h8888;
    LUT4 i1_4_lut_adj_891 (.A(spi_addr_r[6]), .B(n30064), .C(n30155), 
         .D(spi_addr_r[0]), .Z(n26091)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_891.init = 16'h0400;
    LUT4 i1_2_lut_rep_814 (.A(spi_addr_r[6]), .B(spi_addr_r[5]), .Z(n30214)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_814.init = 16'heeee;
    LUT4 i23700_2_lut_3_lut_4_lut (.A(spi_addr_r[6]), .B(spi_addr_r[5]), 
         .C(spi_addr_r[4]), .D(spi_addr_r[1]), .Z(n28402)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23700_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i23780_2_lut_rep_694_3_lut_4_lut (.A(spi_addr_r[6]), .B(spi_addr_r[5]), 
         .C(spi_addr_r[4]), .D(spi_addr_r[7]), .Z(n30094)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23780_2_lut_rep_694_3_lut_4_lut.init = 16'hfffe;
    LUT4 i23784_2_lut_3_lut (.A(spi_addr_r[6]), .B(spi_addr_r[5]), .C(spi_addr_r[7]), 
         .Z(n28486)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i23784_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_892 (.A(n30062), .B(n18440), .C(n26113), .D(n26111), 
         .Z(n26119)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_892.init = 16'hfffd;
    PFUMX i24270 (.BLUT(n29591), .ALUT(n29590), .C0(uart_slot_en[1]), 
          .Z(n29592));
    LUT4 i1_2_lut_adj_893 (.A(spi_addr_r[0]), .B(spi_addr_r[2]), .Z(n26111)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_893.init = 16'heeee;
    LUT4 i3_4_lut (.A(uart_slot_en[0]), .B(n30095), .C(uart_slot_en[3]), 
         .D(pin_io_out_25), .Z(n24734)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 n23552_bdd_3_lut_24363_4_lut (.A(mode_adj_657), .B(n30043), .C(uart_slot_en[0]), 
         .D(n4), .Z(n29590)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam n23552_bdd_3_lut_24363_4_lut.init = 16'hf0e0;
    LUT4 RESET_N_5489_bdd_4_lut (.A(uart_slot_en[2]), .B(pin_io_out_6), 
         .C(n52), .D(mode_adj_658), .Z(n29482)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam RESET_N_5489_bdd_4_lut.init = 16'ha8a0;
    LUT4 i1_3_lut_4_lut (.A(mode_adj_657), .B(n30043), .C(mode_adj_659), 
         .D(pin_io_out_5), .Z(n52)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hfe00;
    LUT4 i1_2_lut_rep_720 (.A(uart_slot_en[1]), .B(uart_slot_en[0]), .Z(n30120)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_720.init = 16'h8888;
    LUT4 i2_2_lut_3_lut (.A(uart_slot_en[1]), .B(uart_slot_en[0]), .C(uart_slot_en[2]), 
         .Z(n23409)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_722 (.A(uart_slot_en[3]), .B(mode_adj_656), .Z(n30122)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_rep_722.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_4_lut_adj_894 (.A(\spi_cmd_r[0] ), .B(spi_addr_r[1]), 
         .C(n28358), .D(\spi_cmd_r[2] ), .Z(n26089)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_894.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_895 (.A(\spi_cmd_r[0] ), .B(spi_addr_r[1]), 
         .C(n25739), .D(\spi_cmd_r[2] ), .Z(n25741)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_895.init = 16'h0080;
    
endmodule
//
// Verilog Description of module \intrpt_ctrl(DEV_ID=4) 
//

module \intrpt_ctrl(DEV_ID=4)  (clk, n30185, \pin_intrpt[12] , intrpt_out_c_4, 
            intrpt_out_N_2926, n31069, \spi_data_out_r_39__N_2863[0] , 
            clear_intrpt, clear_intrpt_N_2930, \spi_data_out_r_39__N_2863[2] , 
            \pin_intrpt[14] , \spi_data_out_r_39__N_2863[1] , \pin_intrpt[13] ) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input n30185;
    input \pin_intrpt[12] ;
    output intrpt_out_c_4;
    input intrpt_out_N_2926;
    input n31069;
    output \spi_data_out_r_39__N_2863[0] ;
    output clear_intrpt;
    input clear_intrpt_N_2930;
    output \spi_data_out_r_39__N_2863[2] ;
    input \pin_intrpt[14] ;
    output \spi_data_out_r_39__N_2863[1] ;
    input \pin_intrpt[13] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire \pin_intrpt[14]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[14] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    wire [2:0]intrpt_in_reg;   // c:/s_links/sources/intrpt_ctrl.v(38[35:48])
    
    wire assert_intrpt;
    wire [2:0]intrpt_in_dly;   // c:/s_links/sources/intrpt_ctrl.v(39[36:49])
    
    wire intrpt_all_edges;
    wire [2:0]intrpt_edge;   // c:/s_links/sources/intrpt_ctrl.v(40[36:47])
    
    FD1S3IX intrpt_in_reg__i0 (.D(\pin_intrpt[12] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i0.GSR = "DISABLED";
    FD1P3IX intrpt_out_359 (.D(n31069), .SP(assert_intrpt), .CD(intrpt_out_N_2926), 
            .CK(clk), .Q(intrpt_out_c_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(92[8] 99[4])
    defparam intrpt_out_359.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i0 (.D(intrpt_in_reg[0]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\pin_intrpt[12] ), .CK(clk), .Q(\spi_data_out_r_39__N_2863[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3IX clear_intrpt_317 (.D(clear_intrpt_N_2930), .CK(clk), .CD(n30185), 
            .Q(clear_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam clear_intrpt_317.GSR = "DISABLED";
    FD1S3IX assert_intrpt_316 (.D(intrpt_all_edges), .CK(clk), .CD(n30185), 
            .Q(assert_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(63[8] 73[4])
    defparam assert_intrpt_316.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\pin_intrpt[14] ), .CK(clk), .Q(\spi_data_out_r_39__N_2863[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\pin_intrpt[13] ), .CK(clk), .Q(\spi_data_out_r_39__N_2863[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i2 (.D(intrpt_in_reg[2]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i1 (.D(intrpt_in_reg[1]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i2 (.D(\pin_intrpt[14] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i1 (.D(\pin_intrpt[13] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i1.GSR = "DISABLED";
    LUT4 i2_4_lut (.A(intrpt_edge[2]), .B(intrpt_in_dly[0]), .C(intrpt_edge[1]), 
         .D(intrpt_in_reg[0]), .Z(intrpt_all_edges)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C+(D)))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i2_4_lut.init = 16'hfbfe;
    LUT4 i1443_2_lut (.A(intrpt_in_dly[2]), .B(intrpt_in_reg[2]), .Z(intrpt_edge[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(46[22:89])
    defparam i1443_2_lut.init = 16'h6666;
    LUT4 i1444_2_lut (.A(intrpt_in_dly[1]), .B(intrpt_in_reg[1]), .Z(intrpt_edge[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(46[22:89])
    defparam i1444_2_lut.init = 16'h6666;
    
endmodule
//
// Verilog Description of module \intrpt_ctrl(DEV_ID=6) 
//

module \intrpt_ctrl(DEV_ID=6)  (clk, n30185, \spi_data_out_r_39__N_3005[0] , 
            \pin_intrpt[18] , intrpt_out_c_6, intrpt_out_N_3068, n31069, 
            \spi_data_out_r_39__N_3005[2] , \pin_intrpt[20] , \spi_data_out_r_39__N_3005[1] , 
            \pin_intrpt[19] , clear_intrpt, clear_intrpt_N_3072) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input n30185;
    output \spi_data_out_r_39__N_3005[0] ;
    input \pin_intrpt[18] ;
    output intrpt_out_c_6;
    input intrpt_out_N_3068;
    input n31069;
    output \spi_data_out_r_39__N_3005[2] ;
    input \pin_intrpt[20] ;
    output \spi_data_out_r_39__N_3005[1] ;
    input \pin_intrpt[19] ;
    output clear_intrpt;
    input clear_intrpt_N_3072;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire \pin_intrpt[20]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[20] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    wire [2:0]intrpt_in_dly;   // c:/s_links/sources/intrpt_ctrl.v(39[36:49])
    wire [2:0]intrpt_in_reg;   // c:/s_links/sources/intrpt_ctrl.v(38[35:48])
    
    wire assert_intrpt, intrpt_all_edges;
    wire [2:0]intrpt_edge;   // c:/s_links/sources/intrpt_ctrl.v(40[36:47])
    
    FD1S3IX intrpt_in_dly__i0 (.D(intrpt_in_reg[0]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\pin_intrpt[18] ), .CK(clk), .Q(\spi_data_out_r_39__N_3005[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1P3IX intrpt_out_359 (.D(n31069), .SP(assert_intrpt), .CD(intrpt_out_N_3068), 
            .CK(clk), .Q(intrpt_out_c_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(92[8] 99[4])
    defparam intrpt_out_359.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i0 (.D(\pin_intrpt[18] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\pin_intrpt[20] ), .CK(clk), .Q(\spi_data_out_r_39__N_3005[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\pin_intrpt[19] ), .CK(clk), .Q(\spi_data_out_r_39__N_3005[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX clear_intrpt_317 (.D(clear_intrpt_N_3072), .CK(clk), .CD(n30185), 
            .Q(clear_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam clear_intrpt_317.GSR = "DISABLED";
    FD1S3IX assert_intrpt_316 (.D(intrpt_all_edges), .CK(clk), .CD(n30185), 
            .Q(assert_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(63[8] 73[4])
    defparam assert_intrpt_316.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i2 (.D(intrpt_in_reg[2]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i1 (.D(intrpt_in_reg[1]), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_dly[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i1 (.D(\pin_intrpt[19] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i2 (.D(\pin_intrpt[20] ), .CK(clk), .CD(n30185), 
            .Q(intrpt_in_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=294, LSE_RLINE=315 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i2.GSR = "DISABLED";
    LUT4 i2_4_lut (.A(intrpt_edge[2]), .B(intrpt_in_dly[0]), .C(intrpt_edge[1]), 
         .D(intrpt_in_reg[0]), .Z(intrpt_all_edges)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C+(D)))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i2_4_lut.init = 16'hfbfe;
    LUT4 i1438_2_lut (.A(intrpt_in_dly[2]), .B(intrpt_in_reg[2]), .Z(intrpt_edge[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(46[22:89])
    defparam i1438_2_lut.init = 16'h6666;
    LUT4 i1439_2_lut (.A(intrpt_in_dly[1]), .B(intrpt_in_reg[1]), .Z(intrpt_edge[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(46[22:89])
    defparam i1439_2_lut.init = 16'h6666;
    
endmodule
//
// Verilog Description of module \status_led(DEV_ID=9) 
//

module \status_led(DEV_ID=9)  (clk, clk_enable_595, n30185, \spi_data_r[0] , 
            \spi_data_out_r_39__N_770[0] , GND_net, n30039, n12435, 
            spi_data_out_r_39__N_810, n12467, \status_cntr[11] , \status_cntr[12] , 
            n18654, EM_STOP, led_sw_c, clk_enable_227, n25212, n4, 
            \spi_data_r[11] , \spi_data_r[10] , \spi_data_r[9] , \spi_data_r[8] , 
            \spi_data_r[7] , \spi_data_r[6] , \spi_data_r[5] , \spi_data_r[4] , 
            \spi_data_r[3] , \spi_data_r[2] , \spi_data_r[1] , pwm, 
            resetn_c, n28562, n57, n6651, pwm_duty_3, n21, n19, 
            n20, n6649, pwm_N_898, n22554, pwm_N_896, n6747, pwm_duty_1, 
            n30020, n20647, n6590, pwm_duty_2, n30102, n29997, \spi_cmd[2] , 
            n27095) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input clk_enable_595;
    input n30185;
    input \spi_data_r[0] ;
    output \spi_data_out_r_39__N_770[0] ;
    input GND_net;
    input n30039;
    input n12435;
    output spi_data_out_r_39__N_810;
    output n12467;
    output \status_cntr[11] ;
    output \status_cntr[12] ;
    output n18654;
    output EM_STOP;
    output led_sw_c;
    input clk_enable_227;
    input n25212;
    output n4;
    input \spi_data_r[11] ;
    input \spi_data_r[10] ;
    input \spi_data_r[9] ;
    input \spi_data_r[8] ;
    input \spi_data_r[7] ;
    input \spi_data_r[6] ;
    input \spi_data_r[5] ;
    input \spi_data_r[4] ;
    input \spi_data_r[3] ;
    input \spi_data_r[2] ;
    input \spi_data_r[1] ;
    output pwm;
    input resetn_c;
    input n28562;
    input n57;
    output n6651;
    input [11:0]pwm_duty_3;
    input n21;
    input n19;
    input n20;
    output n6649;
    output pwm_N_898;
    output n22554;
    output pwm_N_896;
    output n6747;
    input [11:0]pwm_duty_1;
    input n30020;
    input n20647;
    output n6590;
    input [11:0]pwm_duty_2;
    input n30102;
    input n29997;
    input \spi_cmd[2] ;
    input n27095;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire [11:0]pwm_duty;   // c:/s_links/sources/status_led.v(35[30:38])
    
    wire em_stop_flag;
    wire [12:0]pwm_N_899;
    
    wire n21770, n12166;
    wire [12:0]status_cntr;   // c:/s_links/sources/status_led.v(37[32:43])
    
    wire clk_enable_927;
    wire [12:0]n827;
    
    wire n21837, n21838, em_stop_flag_N_917, n28332, n28334, n26277, 
        n26279;
    wire [11:0]pwm_freq_cntr;   // c:/s_links/sources/status_led.v(36[30:43])
    
    wire n21834, n21835, n21839, n21836, n30178, n82, pwm_out_N_893, 
        n12670;
    wire [12:0]n141;
    
    wire n21_c, n19_c, n20_c, n21771, n21773, n22039, n22038, 
        n22037, n22036, n22035, n22034, n21772, n30053, n21_adj_7369, 
        n19_adj_7370, n20_adj_7371, n21_adj_7372, n19_adj_7373, n20_adj_7374;
    wire [11:0]n53;
    
    wire n22138, n22137, n22136, n22135, n22134, n22133, n21_adj_7376, 
        n19_adj_7377, n20_adj_7378;
    
    FD1P3IX pwm_duty__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_595), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(em_stop_flag), .CK(clk), .Q(\spi_data_out_r_39__N_770[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(97[8] 111[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    CCU2D equal_10_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_N_899[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n21770));   // c:/s_links/sources/status_led.v(66[12:41])
    defparam equal_10_0.INIT0 = 16'hF000;
    defparam equal_10_0.INIT1 = 16'h5555;
    defparam equal_10_0.INJECT1_0 = "NO";
    defparam equal_10_0.INJECT1_1 = "YES";
    FD1S3JX em_stop_flag_383 (.D(n12166), .CK(clk), .PD(n30039), .Q(em_stop_flag)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(97[8] 111[4])
    defparam em_stop_flag_383.GSR = "DISABLED";
    FD1P3IX status_cntr_i0_i0 (.D(n827[0]), .SP(clk_enable_927), .CD(n12435), 
            .CK(clk), .Q(status_cntr[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i0.GSR = "DISABLED";
    CCU2D add_395_9 (.A0(status_cntr[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(status_cntr[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21837), .COUT(n21838), .S0(n827[7]), .S1(n827[8]));   // c:/s_links/sources/status_led.v(59[19:34])
    defparam add_395_9.INIT0 = 16'h5aaa;
    defparam add_395_9.INIT1 = 16'h5aaa;
    defparam add_395_9.INJECT1_0 = "NO";
    defparam add_395_9.INJECT1_1 = "NO";
    FD1S3IX i60_343 (.D(em_stop_flag_N_917), .CK(clk), .CD(n30039), .Q(spi_data_out_r_39__N_810)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(97[8] 111[4])
    defparam i60_343.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(n28332), .B(n28334), .C(n26277), .D(n26279), .Z(n12467)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut.init = 16'h1000;
    LUT4 i23630_2_lut (.A(pwm_freq_cntr[2]), .B(pwm_freq_cntr[4]), .Z(n28332)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23630_2_lut.init = 16'heeee;
    LUT4 i23632_2_lut (.A(pwm_freq_cntr[11]), .B(pwm_freq_cntr[7]), .Z(n28334)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23632_2_lut.init = 16'heeee;
    CCU2D add_395_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(status_cntr[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n21834), .S1(n827[0]));   // c:/s_links/sources/status_led.v(59[19:34])
    defparam add_395_1.INIT0 = 16'hF000;
    defparam add_395_1.INIT1 = 16'h5555;
    defparam add_395_1.INJECT1_0 = "NO";
    defparam add_395_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_866 (.A(pwm_freq_cntr[8]), .B(pwm_freq_cntr[3]), .C(pwm_freq_cntr[10]), 
         .D(pwm_freq_cntr[6]), .Z(n26277)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_866.init = 16'h8000;
    CCU2D add_395_3 (.A0(status_cntr[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(status_cntr[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21834), .COUT(n21835), .S0(n827[1]), .S1(n827[2]));   // c:/s_links/sources/status_led.v(59[19:34])
    defparam add_395_3.INIT0 = 16'h5aaa;
    defparam add_395_3.INIT1 = 16'h5aaa;
    defparam add_395_3.INJECT1_0 = "NO";
    defparam add_395_3.INJECT1_1 = "NO";
    CCU2D add_395_13 (.A0(\status_cntr[11] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\status_cntr[12] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21839), .S0(n827[11]), .S1(n827[12]));   // c:/s_links/sources/status_led.v(59[19:34])
    defparam add_395_13.INIT0 = 16'h5aaa;
    defparam add_395_13.INIT1 = 16'h5aaa;
    defparam add_395_13.INJECT1_0 = "NO";
    defparam add_395_13.INJECT1_1 = "NO";
    CCU2D add_395_7 (.A0(status_cntr[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(status_cntr[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21836), .COUT(n21837), .S0(n827[5]), .S1(n827[6]));   // c:/s_links/sources/status_led.v(59[19:34])
    defparam add_395_7.INIT0 = 16'h5aaa;
    defparam add_395_7.INIT1 = 16'h5aaa;
    defparam add_395_7.INJECT1_0 = "NO";
    defparam add_395_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_867 (.A(pwm_freq_cntr[1]), .B(pwm_freq_cntr[0]), .C(pwm_freq_cntr[9]), 
         .D(pwm_freq_cntr[5]), .Z(n26279)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_867.init = 16'h8000;
    LUT4 i1_4_lut_adj_868 (.A(\status_cntr[11] ), .B(\status_cntr[12] ), 
         .C(n30178), .D(n82), .Z(n18654)) /* synthesis lut_function=(A (B)+!A (B (C (D)))) */ ;   // c:/s_links/sources/status_led.v(37[32:43])
    defparam i1_4_lut_adj_868.init = 16'hc888;
    LUT4 i1_4_lut_adj_869 (.A(status_cntr[5]), .B(status_cntr[7]), .C(status_cntr[6]), 
         .D(status_cntr[4]), .Z(n82)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;   // c:/s_links/sources/status_led.v(37[32:43])
    defparam i1_4_lut_adj_869.init = 16'heccc;
    FD1S3IX EM_STOP_338 (.D(pwm_out_N_893), .CK(clk), .CD(n30185), .Q(EM_STOP)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam EM_STOP_338.GSR = "DISABLED";
    FD1P3AX pwm_out_337 (.D(n25212), .SP(clk_enable_227), .CK(clk), .Q(led_sw_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_out_337.GSR = "DISABLED";
    LUT4 i4_3_lut_4_lut (.A(status_cntr[7]), .B(n30178), .C(status_cntr[5]), 
         .D(status_cntr[6]), .Z(n4)) /* synthesis lut_function=(!(A (B (C+(D))))) */ ;   // c:/s_links/sources/status_led.v(37[32:43])
    defparam i4_3_lut_4_lut.init = 16'h777f;
    LUT4 i7804_2_lut (.A(em_stop_flag_N_917), .B(em_stop_flag), .Z(n12166)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/s_links/sources/status_led.v(97[8] 111[4])
    defparam i7804_2_lut.init = 16'h4444;
    CCU2D add_395_5 (.A0(status_cntr[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(status_cntr[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21835), .COUT(n21836), .S0(n827[3]), .S1(n827[4]));   // c:/s_links/sources/status_led.v(59[19:34])
    defparam add_395_5.INIT0 = 16'h5aaa;
    defparam add_395_5.INIT1 = 16'h5aaa;
    defparam add_395_5.INJECT1_0 = "NO";
    defparam add_395_5.INJECT1_1 = "NO";
    CCU2D add_395_11 (.A0(status_cntr[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(status_cntr[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21838), .COUT(n21839), .S0(n827[9]), .S1(n827[10]));   // c:/s_links/sources/status_led.v(59[19:34])
    defparam add_395_11.INIT0 = 16'h5aaa;
    defparam add_395_11.INIT1 = 16'h5aaa;
    defparam add_395_11.INJECT1_0 = "NO";
    defparam add_395_11.INJECT1_1 = "NO";
    FD1P3IX pwm_duty__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_595), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i11.GSR = "DISABLED";
    FD1P3IX pwm_duty__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_595), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i10.GSR = "DISABLED";
    FD1P3IX pwm_duty__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_595), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i9.GSR = "DISABLED";
    FD1P3IX pwm_duty__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_595), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i8.GSR = "DISABLED";
    FD1P3IX pwm_duty__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_595), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i7.GSR = "DISABLED";
    FD1P3IX pwm_duty__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_595), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i6.GSR = "DISABLED";
    FD1P3IX pwm_duty__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_595), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i5.GSR = "DISABLED";
    FD1P3IX pwm_duty__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_595), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i4.GSR = "DISABLED";
    FD1P3IX pwm_duty__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_595), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i3.GSR = "DISABLED";
    FD1P3IX pwm_duty__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_595), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i2.GSR = "DISABLED";
    FD1P3IX pwm_duty__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_595), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i1.GSR = "DISABLED";
    FD1P3AX pwm_341 (.D(n28562), .SP(resetn_c), .CK(clk), .Q(pwm)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_341.GSR = "DISABLED";
    LUT4 i8106_2_lut (.A(resetn_c), .B(n12467), .Z(n12670)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam i8106_2_lut.init = 16'h8888;
    LUT4 i1_2_lut (.A(n12467), .B(n827[4]), .Z(n141[4])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_870 (.A(n12467), .B(n827[8]), .Z(n141[8])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_870.init = 16'h8888;
    LUT4 i1_2_lut_adj_871 (.A(n12467), .B(n827[9]), .Z(n141[9])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_871.init = 16'h8888;
    LUT4 i1_2_lut_adj_872 (.A(n12467), .B(n827[6]), .Z(n141[6])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_872.init = 16'h8888;
    LUT4 i1_2_lut_adj_873 (.A(n12467), .B(n827[7]), .Z(n141[7])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_873.init = 16'h8888;
    LUT4 i1_2_lut_adj_874 (.A(n12467), .B(n827[10]), .Z(n141[10])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_874.init = 16'h8888;
    LUT4 i1_4_lut_adj_875 (.A(n21_c), .B(n57), .C(n19_c), .D(n20_c), 
         .Z(n6651)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // c:/s_links/sources/status_led.v(98[6:24])
    defparam i1_4_lut_adj_875.init = 16'h3332;
    LUT4 i9_4_lut (.A(pwm_duty_3[3]), .B(pwm_duty_3[0]), .C(pwm_duty_3[8]), 
         .D(pwm_duty_3[2]), .Z(n21_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(57[38:48])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i7_4_lut (.A(pwm_duty_3[6]), .B(pwm_duty_3[5]), .C(pwm_duty_3[4]), 
         .D(pwm_duty_3[7]), .Z(n19_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(57[38:48])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i8_4_lut (.A(pwm_duty_3[9]), .B(pwm_duty_3[1]), .C(pwm_duty_3[10]), 
         .D(pwm_duty_3[11]), .Z(n20_c)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(57[38:48])
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_876 (.A(n21), .B(n57), .C(n19), .D(n20), .Z(n6649)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // c:/s_links/sources/status_led.v(98[6:24])
    defparam i1_4_lut_adj_876.init = 16'h3332;
    CCU2D equal_10_9 (.A0(pwm_N_899[11]), .B0(pwm_freq_cntr[11]), .C0(pwm_N_899[10]), 
          .D0(pwm_freq_cntr[10]), .A1(pwm_N_899[9]), .B1(pwm_freq_cntr[9]), 
          .C1(pwm_N_899[8]), .D1(pwm_freq_cntr[8]), .CIN(n21770), .COUT(n21771));
    defparam equal_10_9.INIT0 = 16'h9009;
    defparam equal_10_9.INIT1 = 16'h9009;
    defparam equal_10_9.INJECT1_0 = "YES";
    defparam equal_10_9.INJECT1_1 = "YES";
    CCU2D equal_10_13 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21773), 
          .S0(pwm_N_898));
    defparam equal_10_13.INIT0 = 16'hFFFF;
    defparam equal_10_13.INIT1 = 16'h0000;
    defparam equal_10_13.INJECT1_0 = "NO";
    defparam equal_10_13.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_13 (.A0(pwm_duty[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n22039), .S0(pwm_N_899[11]), .S1(pwm_N_899[12]));   // c:/s_links/sources/status_led.v(66[29:41])
    defparam sub_14_add_2_13.INIT0 = 16'h5555;
    defparam sub_14_add_2_13.INIT1 = 16'hffff;
    defparam sub_14_add_2_13.INJECT1_0 = "NO";
    defparam sub_14_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_11 (.A0(pwm_duty[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22038), .COUT(n22039), .S0(pwm_N_899[9]), 
          .S1(pwm_N_899[10]));   // c:/s_links/sources/status_led.v(66[29:41])
    defparam sub_14_add_2_11.INIT0 = 16'h5555;
    defparam sub_14_add_2_11.INIT1 = 16'h5555;
    defparam sub_14_add_2_11.INJECT1_0 = "NO";
    defparam sub_14_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_9 (.A0(pwm_duty[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22037), .COUT(n22038), .S0(pwm_N_899[7]), 
          .S1(pwm_N_899[8]));   // c:/s_links/sources/status_led.v(66[29:41])
    defparam sub_14_add_2_9.INIT0 = 16'h5555;
    defparam sub_14_add_2_9.INIT1 = 16'h5555;
    defparam sub_14_add_2_9.INJECT1_0 = "NO";
    defparam sub_14_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_7 (.A0(pwm_duty[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22036), .COUT(n22037), .S0(pwm_N_899[5]), 
          .S1(pwm_N_899[6]));   // c:/s_links/sources/status_led.v(66[29:41])
    defparam sub_14_add_2_7.INIT0 = 16'h5555;
    defparam sub_14_add_2_7.INIT1 = 16'h5555;
    defparam sub_14_add_2_7.INJECT1_0 = "NO";
    defparam sub_14_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_5 (.A0(pwm_duty[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22035), .COUT(n22036), .S0(pwm_N_899[3]), 
          .S1(pwm_N_899[4]));   // c:/s_links/sources/status_led.v(66[29:41])
    defparam sub_14_add_2_5.INIT0 = 16'h5555;
    defparam sub_14_add_2_5.INIT1 = 16'h5555;
    defparam sub_14_add_2_5.INJECT1_0 = "NO";
    defparam sub_14_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_3 (.A0(pwm_duty[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22034), .COUT(n22035), .S0(pwm_N_899[1]), 
          .S1(pwm_N_899[2]));   // c:/s_links/sources/status_led.v(66[29:41])
    defparam sub_14_add_2_3.INIT0 = 16'h5555;
    defparam sub_14_add_2_3.INIT1 = 16'h5555;
    defparam sub_14_add_2_3.INJECT1_0 = "NO";
    defparam sub_14_add_2_3.INJECT1_1 = "NO";
    CCU2D equal_10_13_17464 (.A0(pwm_N_899[3]), .B0(pwm_freq_cntr[3]), .C0(pwm_N_899[2]), 
          .D0(pwm_freq_cntr[2]), .A1(pwm_N_899[1]), .B1(pwm_freq_cntr[1]), 
          .C1(pwm_N_899[0]), .D1(pwm_freq_cntr[0]), .CIN(n21772), .COUT(n21773));
    defparam equal_10_13_17464.INIT0 = 16'h9009;
    defparam equal_10_13_17464.INIT1 = 16'h9009;
    defparam equal_10_13_17464.INJECT1_0 = "YES";
    defparam equal_10_13_17464.INJECT1_1 = "YES";
    CCU2D sub_14_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_duty[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n22034), .S1(pwm_N_899[0]));   // c:/s_links/sources/status_led.v(66[29:41])
    defparam sub_14_add_2_1.INIT0 = 16'hF000;
    defparam sub_14_add_2_1.INIT1 = 16'h5555;
    defparam sub_14_add_2_1.INJECT1_0 = "NO";
    defparam sub_14_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_3_lut (.A(\status_cntr[12] ), .B(n22554), .C(\status_cntr[11] ), 
         .Z(pwm_out_N_893)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_877 (.A(status_cntr[5]), .B(n30053), .C(status_cntr[6]), 
         .D(status_cntr[4]), .Z(n22554)) /* synthesis lut_function=(A (B (C))+!A (B (C (D)))) */ ;   // c:/s_links/sources/status_led.v(37[32:43])
    defparam i1_4_lut_adj_877.init = 16'hc080;
    CCU2D equal_10_11 (.A0(pwm_N_899[7]), .B0(pwm_freq_cntr[7]), .C0(pwm_N_899[6]), 
          .D0(pwm_freq_cntr[6]), .A1(pwm_N_899[5]), .B1(pwm_freq_cntr[5]), 
          .C1(pwm_N_899[4]), .D1(pwm_freq_cntr[4]), .CIN(n21771), .COUT(n21772));
    defparam equal_10_11.INIT0 = 16'h9009;
    defparam equal_10_11.INIT1 = 16'h9009;
    defparam equal_10_11.INJECT1_0 = "YES";
    defparam equal_10_11.INJECT1_1 = "YES";
    LUT4 i1_4_lut_adj_878 (.A(n12467), .B(n21_adj_7369), .C(n19_adj_7370), 
         .D(n20_adj_7371), .Z(pwm_N_896)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_878.init = 16'haaa8;
    LUT4 i9_4_lut_adj_879 (.A(pwm_duty[11]), .B(pwm_duty[8]), .C(pwm_duty[3]), 
         .D(pwm_duty[0]), .Z(n21_adj_7369)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/status_led.v(61[8:23])
    defparam i9_4_lut_adj_879.init = 16'hfffe;
    LUT4 i7_4_lut_adj_880 (.A(pwm_duty[4]), .B(pwm_duty[9]), .C(pwm_duty[10]), 
         .D(pwm_duty[1]), .Z(n19_adj_7370)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/status_led.v(61[8:23])
    defparam i7_4_lut_adj_880.init = 16'hfffe;
    LUT4 i8_4_lut_adj_881 (.A(pwm_duty[6]), .B(pwm_duty[2]), .C(pwm_duty[5]), 
         .D(pwm_duty[7]), .Z(n20_adj_7371)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/status_led.v(61[8:23])
    defparam i8_4_lut_adj_881.init = 16'hfffe;
    LUT4 i1_3_lut_rep_778 (.A(status_cntr[8]), .B(status_cntr[9]), .C(status_cntr[10]), 
         .Z(n30178)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam i1_3_lut_rep_778.init = 16'h8080;
    LUT4 i1_2_lut_rep_653_4_lut (.A(status_cntr[8]), .B(status_cntr[9]), 
         .C(status_cntr[10]), .D(status_cntr[7]), .Z(n30053)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam i1_2_lut_rep_653_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_882 (.A(n21_adj_7372), .B(n57), .C(n19_adj_7373), 
         .D(n20_adj_7374), .Z(n6747)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // c:/s_links/sources/status_led.v(98[6:24])
    defparam i1_4_lut_adj_882.init = 16'h3332;
    LUT4 i9_4_lut_adj_883 (.A(pwm_duty_1[5]), .B(pwm_duty_1[10]), .C(pwm_duty_1[6]), 
         .D(pwm_duty_1[2]), .Z(n21_adj_7372)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(55[38:48])
    defparam i9_4_lut_adj_883.init = 16'hfffe;
    LUT4 i7_4_lut_adj_884 (.A(pwm_duty_1[8]), .B(pwm_duty_1[3]), .C(pwm_duty_1[4]), 
         .D(pwm_duty_1[7]), .Z(n19_adj_7373)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(55[38:48])
    defparam i7_4_lut_adj_884.init = 16'hfffe;
    LUT4 i8_4_lut_adj_885 (.A(pwm_duty_1[9]), .B(pwm_duty_1[11]), .C(pwm_duty_1[0]), 
         .D(pwm_duty_1[1]), .Z(n20_adj_7374)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(55[38:48])
    defparam i8_4_lut_adj_885.init = 16'hfffe;
    FD1P3IX pwm_freq_cntr_1776__i11 (.D(n53[11]), .SP(resetn_c), .CD(n12670), 
            .CK(clk), .Q(pwm_freq_cntr[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776__i11.GSR = "DISABLED";
    CCU2D pwm_freq_cntr_1776_add_4_13 (.A0(pwm_freq_cntr[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22138), .S0(n53[11]));   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776_add_4_13.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1776_add_4_13.INIT1 = 16'h0000;
    defparam pwm_freq_cntr_1776_add_4_13.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1776_add_4_13.INJECT1_1 = "NO";
    FD1P3IX pwm_freq_cntr_1776__i1 (.D(n53[1]), .SP(resetn_c), .CD(n12670), 
            .CK(clk), .Q(pwm_freq_cntr[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776__i1.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_1776__i5 (.D(n53[5]), .SP(resetn_c), .CD(n12670), 
            .CK(clk), .Q(pwm_freq_cntr[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776__i5.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_1776__i8 (.D(n53[8]), .SP(resetn_c), .CD(n12670), 
            .CK(clk), .Q(pwm_freq_cntr[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776__i8.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_1776__i2 (.D(n53[2]), .SP(resetn_c), .CD(n12670), 
            .CK(clk), .Q(pwm_freq_cntr[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776__i2.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_1776__i6 (.D(n53[6]), .SP(resetn_c), .CD(n12670), 
            .CK(clk), .Q(pwm_freq_cntr[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776__i6.GSR = "DISABLED";
    CCU2D pwm_freq_cntr_1776_add_4_11 (.A0(pwm_freq_cntr[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n22137), .COUT(n22138), .S0(n53[9]), 
          .S1(n53[10]));   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776_add_4_11.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1776_add_4_11.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1776_add_4_11.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1776_add_4_11.INJECT1_1 = "NO";
    FD1P3IX pwm_freq_cntr_1776__i9 (.D(n53[9]), .SP(resetn_c), .CD(n12670), 
            .CK(clk), .Q(pwm_freq_cntr[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776__i9.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_1776__i3 (.D(n53[3]), .SP(resetn_c), .CD(n12670), 
            .CK(clk), .Q(pwm_freq_cntr[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776__i3.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_1776__i4 (.D(n53[4]), .SP(resetn_c), .CD(n12670), 
            .CK(clk), .Q(pwm_freq_cntr[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776__i4.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_1776__i7 (.D(n53[7]), .SP(resetn_c), .CD(n12670), 
            .CK(clk), .Q(pwm_freq_cntr[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776__i7.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_1776__i10 (.D(n53[10]), .SP(resetn_c), .CD(n12670), 
            .CK(clk), .Q(pwm_freq_cntr[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776__i10.GSR = "DISABLED";
    FD1P3JX status_cntr_i0_i4 (.D(n141[4]), .SP(clk_enable_927), .PD(n30020), 
            .CK(clk), .Q(status_cntr[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i4.GSR = "DISABLED";
    FD1P3JX status_cntr_i0_i8 (.D(n141[8]), .SP(clk_enable_927), .PD(n30020), 
            .CK(clk), .Q(status_cntr[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i8.GSR = "DISABLED";
    FD1P3IX status_cntr_i0_i11 (.D(n827[11]), .SP(clk_enable_927), .CD(n12435), 
            .CK(clk), .Q(\status_cntr[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i11.GSR = "DISABLED";
    FD1P3IX status_cntr_i0_i5 (.D(n827[5]), .SP(clk_enable_927), .CD(n12435), 
            .CK(clk), .Q(status_cntr[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i5.GSR = "DISABLED";
    FD1P3JX status_cntr_i0_i9 (.D(n141[9]), .SP(clk_enable_927), .PD(n30020), 
            .CK(clk), .Q(status_cntr[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i9.GSR = "DISABLED";
    FD1P3IX status_cntr_i0_i12 (.D(n827[12]), .SP(clk_enable_927), .CD(n12435), 
            .CK(clk), .Q(\status_cntr[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i12.GSR = "DISABLED";
    FD1P3IX status_cntr_i0_i2 (.D(n827[2]), .SP(clk_enable_927), .CD(n12435), 
            .CK(clk), .Q(status_cntr[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i2.GSR = "DISABLED";
    FD1P3JX status_cntr_i0_i6 (.D(n141[6]), .SP(clk_enable_927), .PD(n30020), 
            .CK(clk), .Q(status_cntr[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i6.GSR = "DISABLED";
    FD1P3IX status_cntr_i0_i3 (.D(n827[3]), .SP(clk_enable_927), .CD(n12435), 
            .CK(clk), .Q(status_cntr[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i3.GSR = "DISABLED";
    FD1P3JX status_cntr_i0_i7 (.D(n141[7]), .SP(clk_enable_927), .PD(n30020), 
            .CK(clk), .Q(status_cntr[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i7.GSR = "DISABLED";
    FD1P3JX status_cntr_i0_i10 (.D(n141[10]), .SP(clk_enable_927), .PD(n30020), 
            .CK(clk), .Q(status_cntr[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i10.GSR = "DISABLED";
    CCU2D pwm_freq_cntr_1776_add_4_9 (.A0(pwm_freq_cntr[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n22136), .COUT(n22137), .S0(n53[7]), 
          .S1(n53[8]));   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776_add_4_9.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1776_add_4_9.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1776_add_4_9.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1776_add_4_9.INJECT1_1 = "NO";
    FD1P3IX status_cntr_i0_i1 (.D(n827[1]), .SP(clk_enable_927), .CD(n12435), 
            .CK(clk), .Q(status_cntr[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=219, LSE_RLINE=236 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i1.GSR = "DISABLED";
    CCU2D pwm_freq_cntr_1776_add_4_7 (.A0(pwm_freq_cntr[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n22135), .COUT(n22136), .S0(n53[5]), 
          .S1(n53[6]));   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776_add_4_7.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1776_add_4_7.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1776_add_4_7.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1776_add_4_7.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1776_add_4_5 (.A0(pwm_freq_cntr[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n22134), .COUT(n22135), .S0(n53[3]), 
          .S1(n53[4]));   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776_add_4_5.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1776_add_4_5.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1776_add_4_5.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1776_add_4_5.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1776_add_4_3 (.A0(pwm_freq_cntr[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n22133), .COUT(n22134), .S0(n53[1]), 
          .S1(n53[2]));   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776_add_4_3.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1776_add_4_3.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1776_add_4_3.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1776_add_4_3.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1776_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_freq_cntr[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n22133), .S1(n53[0]));   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776_add_4_1.INIT0 = 16'hF000;
    defparam pwm_freq_cntr_1776_add_4_1.INIT1 = 16'h0555;
    defparam pwm_freq_cntr_1776_add_4_1.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1776_add_4_1.INJECT1_1 = "NO";
    FD1P3IX pwm_freq_cntr_1776__i0 (.D(n53[0]), .SP(resetn_c), .CD(n12670), 
            .CK(clk), .Q(pwm_freq_cntr[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_1776__i0.GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut (.A(n18654), .B(n20647), .C(n12467), .D(resetn_c), 
         .Z(clk_enable_927)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfe00;
    LUT4 i1_4_lut_adj_886 (.A(n21_adj_7376), .B(n57), .C(n19_adj_7377), 
         .D(n20_adj_7378), .Z(n6590)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // c:/s_links/sources/status_led.v(98[6:24])
    defparam i1_4_lut_adj_886.init = 16'h3332;
    LUT4 i9_4_lut_adj_887 (.A(pwm_duty_2[7]), .B(pwm_duty_2[9]), .C(pwm_duty_2[8]), 
         .D(pwm_duty_2[2]), .Z(n21_adj_7376)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(56[38:48])
    defparam i9_4_lut_adj_887.init = 16'hfffe;
    LUT4 i7_4_lut_adj_888 (.A(pwm_duty_2[11]), .B(pwm_duty_2[5]), .C(pwm_duty_2[4]), 
         .D(pwm_duty_2[6]), .Z(n19_adj_7377)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(56[38:48])
    defparam i7_4_lut_adj_888.init = 16'hfffe;
    LUT4 i8_4_lut_adj_889 (.A(pwm_duty_2[0]), .B(pwm_duty_2[1]), .C(pwm_duty_2[10]), 
         .D(pwm_duty_2[3]), .Z(n20_adj_7378)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(56[38:48])
    defparam i8_4_lut_adj_889.init = 16'hfffe;
    LUT4 i24136_4_lut (.A(n30102), .B(n29997), .C(\spi_cmd[2] ), .D(n27095), 
         .Z(em_stop_flag_N_917)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/s_links/sources/status_led.v(102[15:46])
    defparam i24136_4_lut.init = 16'h0010;
    
endmodule
//
// Verilog Description of module pll
//

module pll (clk_in_c, clk_100k, clk_1MHz, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input clk_in_c;
    output clk_100k;
    output clk_1MHz;
    input GND_net;
    
    wire clk_in_c /* synthesis is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(16[27:33])
    wire clk_100k /* synthesis SET_AS_NETWORK=clk_100k, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(134[6:14])
    wire clk_1MHz /* synthesis SET_AS_NETWORK=clk_1MHz, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(136[6:14])
    
    wire CLKFB_t;
    
    EHXPLLJ PLLInst_0 (.CLKI(clk_in_c), .CLKFB(CLKFB_t), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(GND_net), .PLLRST(GND_net), .PLLSTB(GND_net), 
            .PLLWE(GND_net), .PLLDATI0(GND_net), .PLLDATI1(GND_net), .PLLDATI2(GND_net), 
            .PLLDATI3(GND_net), .PLLDATI4(GND_net), .PLLDATI5(GND_net), 
            .PLLDATI6(GND_net), .PLLDATI7(GND_net), .PLLADDR0(GND_net), 
            .PLLADDR1(GND_net), .PLLADDR2(GND_net), .PLLADDR3(GND_net), 
            .PLLADDR4(GND_net), .CLKOS(clk_100k), .CLKOS3(clk_1MHz), .CLKINTFB(CLKFB_t)) /* synthesis FREQUENCY_PIN_CLKOS3="1.000000", FREQUENCY_PIN_CLKOS2="0.020000", FREQUENCY_PIN_CLKOS="0.100000", FREQUENCY_PIN_CLKOP="96.000000", FREQUENCY_PIN_CLKI="12.000000", ICP_CURRENT="9", LPF_RESISTOR="4", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=100, LSE_LLINE=140, LSE_RLINE=140 */ ;   // c:/s_links/sources/mcm_top.v(140[5:100])
    defparam PLLInst_0.CLKI_DIV = 1;
    defparam PLLInst_0.CLKFB_DIV = 8;
    defparam PLLInst_0.CLKOP_DIV = 3;
    defparam PLLInst_0.CLKOS_DIV = 120;
    defparam PLLInst_0.CLKOS2_DIV = 120;
    defparam PLLInst_0.CLKOS3_DIV = 12;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "ENABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "ENABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "ENABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 2;
    defparam PLLInst_0.CLKOS_CPHASE = 119;
    defparam PLLInst_0.CLKOS2_CPHASE = 119;
    defparam PLLInst_0.CLKOS3_CPHASE = 11;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "INT_DIVA";
    defparam PLLInst_0.FRACN_ENABLE = "DISABLED";
    defparam PLLInst_0.FRACN_DIV = 0;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "DISABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 3;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module pwm_controller
//

module pwm_controller (\pwm_out[0] , clk, clk_enable_15, n2109, clk_enable_263, 
            n30185, \spi_data_r[0] , clk_enable_638, \spi_data_r[11] , 
            \spi_data_r[10] , \spi_data_r[9] , \spi_data_r[8] , \spi_data_r[7] , 
            \spi_data_r[6] , \spi_data_r[5] , \spi_data_r[4] , \spi_data_r[3] , 
            \spi_data_r[2] , \spi_data_r[1] , GND_net, pwm_out_N_3153, 
            pwm_out_N_3169, resetn_c) /* synthesis syn_module_defined=1 */ ;
    output \pwm_out[0] ;
    input clk;
    input clk_enable_15;
    input n2109;
    input clk_enable_263;
    input n30185;
    input \spi_data_r[0] ;
    input clk_enable_638;
    input \spi_data_r[11] ;
    input \spi_data_r[10] ;
    input \spi_data_r[9] ;
    input \spi_data_r[8] ;
    input \spi_data_r[7] ;
    input \spi_data_r[6] ;
    input \spi_data_r[5] ;
    input \spi_data_r[4] ;
    input \spi_data_r[3] ;
    input \spi_data_r[2] ;
    input \spi_data_r[1] ;
    input GND_net;
    output pwm_out_N_3153;
    output pwm_out_N_3169;
    input resetn_c;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    
    wire n25197;
    wire [11:0]pwm_freq_cntr;   // c:/s_links/sources/pwm_controller.v(30[30:43])
    wire [11:0]n53;
    wire [11:0]pwm_freq;   // c:/s_links/sources/pwm_controller.v(28[30:38])
    wire [11:0]pwm_duty;   // c:/s_links/sources/pwm_controller.v(29[30:38])
    
    wire n21866, n21781, n21865, n21864, n21863, n21862, n21780;
    wire [12:0]pwm_out_N_3154;
    wire [12:0]pwm_out_N_3170;
    
    wire n21774, n21861, n21779, n21778, n22032, n22031, n21777, 
        n22030, n22029, n22028, n22027, n22025, n22024, n22023, 
        n22022, n21776, n22021, n22020, n21775, n28249, n28243, 
        n28245, n28231;
    
    FD1P3AX pwm_out_40 (.D(n25197), .SP(clk_enable_15), .CK(clk), .Q(\pwm_out[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(53[8] 75[4])
    defparam pwm_out_40.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1777__i0 (.D(n53[0]), .CK(clk), .CD(n2109), 
            .Q(pwm_freq_cntr[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777__i0.GSR = "DISABLED";
    FD1P3IX pwm_freq__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_263), .CD(n30185), 
            .CK(clk), .Q(pwm_freq[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(34[8] 41[4])
    defparam pwm_freq__i0.GSR = "DISABLED";
    FD1P3IX pwm_duty__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_638), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(43[8] 50[4])
    defparam pwm_duty__i0.GSR = "DISABLED";
    FD1P3IX pwm_freq__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_263), .CD(n30185), 
            .CK(clk), .Q(pwm_freq[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(34[8] 41[4])
    defparam pwm_freq__i11.GSR = "DISABLED";
    FD1P3IX pwm_freq__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_263), .CD(n30185), 
            .CK(clk), .Q(pwm_freq[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(34[8] 41[4])
    defparam pwm_freq__i10.GSR = "DISABLED";
    FD1P3IX pwm_freq__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_263), .CD(n30185), 
            .CK(clk), .Q(pwm_freq[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(34[8] 41[4])
    defparam pwm_freq__i9.GSR = "DISABLED";
    FD1P3IX pwm_freq__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_263), .CD(n30185), 
            .CK(clk), .Q(pwm_freq[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(34[8] 41[4])
    defparam pwm_freq__i8.GSR = "DISABLED";
    FD1P3IX pwm_freq__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_263), .CD(n30185), 
            .CK(clk), .Q(pwm_freq[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(34[8] 41[4])
    defparam pwm_freq__i7.GSR = "DISABLED";
    FD1P3IX pwm_freq__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_263), .CD(n30185), 
            .CK(clk), .Q(pwm_freq[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(34[8] 41[4])
    defparam pwm_freq__i6.GSR = "DISABLED";
    FD1P3IX pwm_freq__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_263), .CD(n30185), 
            .CK(clk), .Q(pwm_freq[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(34[8] 41[4])
    defparam pwm_freq__i5.GSR = "DISABLED";
    FD1P3IX pwm_freq__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_263), .CD(n30185), 
            .CK(clk), .Q(pwm_freq[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(34[8] 41[4])
    defparam pwm_freq__i4.GSR = "DISABLED";
    FD1P3IX pwm_freq__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_263), .CD(n30185), 
            .CK(clk), .Q(pwm_freq[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(34[8] 41[4])
    defparam pwm_freq__i3.GSR = "DISABLED";
    FD1P3IX pwm_freq__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_263), .CD(n30185), 
            .CK(clk), .Q(pwm_freq[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(34[8] 41[4])
    defparam pwm_freq__i2.GSR = "DISABLED";
    FD1P3IX pwm_freq__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_263), .CD(n30185), 
            .CK(clk), .Q(pwm_freq[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(34[8] 41[4])
    defparam pwm_freq__i1.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1777__i11 (.D(n53[11]), .CK(clk), .CD(n2109), 
            .Q(pwm_freq_cntr[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777__i11.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1777__i10 (.D(n53[10]), .CK(clk), .CD(n2109), 
            .Q(pwm_freq_cntr[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777__i10.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1777__i9 (.D(n53[9]), .CK(clk), .CD(n2109), 
            .Q(pwm_freq_cntr[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777__i9.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1777__i8 (.D(n53[8]), .CK(clk), .CD(n2109), 
            .Q(pwm_freq_cntr[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777__i8.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1777__i7 (.D(n53[7]), .CK(clk), .CD(n2109), 
            .Q(pwm_freq_cntr[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777__i7.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1777__i6 (.D(n53[6]), .CK(clk), .CD(n2109), 
            .Q(pwm_freq_cntr[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777__i6.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1777__i5 (.D(n53[5]), .CK(clk), .CD(n2109), 
            .Q(pwm_freq_cntr[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777__i5.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1777__i4 (.D(n53[4]), .CK(clk), .CD(n2109), 
            .Q(pwm_freq_cntr[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777__i4.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1777__i3 (.D(n53[3]), .CK(clk), .CD(n2109), 
            .Q(pwm_freq_cntr[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777__i3.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1777__i2 (.D(n53[2]), .CK(clk), .CD(n2109), 
            .Q(pwm_freq_cntr[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777__i2.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1777__i1 (.D(n53[1]), .CK(clk), .CD(n2109), 
            .Q(pwm_freq_cntr[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777__i1.GSR = "DISABLED";
    FD1P3IX pwm_duty__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_638), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(43[8] 50[4])
    defparam pwm_duty__i1.GSR = "DISABLED";
    FD1P3IX pwm_duty__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_638), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(43[8] 50[4])
    defparam pwm_duty__i2.GSR = "DISABLED";
    FD1P3IX pwm_duty__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_638), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(43[8] 50[4])
    defparam pwm_duty__i3.GSR = "DISABLED";
    FD1P3IX pwm_duty__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_638), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(43[8] 50[4])
    defparam pwm_duty__i4.GSR = "DISABLED";
    FD1P3IX pwm_duty__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_638), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(43[8] 50[4])
    defparam pwm_duty__i5.GSR = "DISABLED";
    FD1P3IX pwm_duty__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_638), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(43[8] 50[4])
    defparam pwm_duty__i6.GSR = "DISABLED";
    FD1P3IX pwm_duty__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_638), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(43[8] 50[4])
    defparam pwm_duty__i7.GSR = "DISABLED";
    FD1P3IX pwm_duty__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_638), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(43[8] 50[4])
    defparam pwm_duty__i8.GSR = "DISABLED";
    FD1P3IX pwm_duty__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_638), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(43[8] 50[4])
    defparam pwm_duty__i9.GSR = "DISABLED";
    FD1P3IX pwm_duty__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_638), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(43[8] 50[4])
    defparam pwm_duty__i10.GSR = "DISABLED";
    FD1P3IX pwm_duty__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_638), .CD(n30185), 
            .CK(clk), .Q(pwm_duty[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=4, LSE_LLINE=327, LSE_RLINE=339 */ ;   // c:/s_links/sources/pwm_controller.v(43[8] 50[4])
    defparam pwm_duty__i11.GSR = "DISABLED";
    CCU2D pwm_freq_cntr_1777_add_4_13 (.A0(pwm_freq_cntr[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21866), .S0(n53[11]));   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777_add_4_13.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1777_add_4_13.INIT1 = 16'h0000;
    defparam pwm_freq_cntr_1777_add_4_13.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1777_add_4_13.INJECT1_1 = "NO";
    CCU2D equal_54_13 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21781), 
          .S0(pwm_out_N_3153));
    defparam equal_54_13.INIT0 = 16'hFFFF;
    defparam equal_54_13.INIT1 = 16'h0000;
    defparam equal_54_13.INJECT1_0 = "NO";
    defparam equal_54_13.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1777_add_4_11 (.A0(pwm_freq_cntr[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n21865), .COUT(n21866), .S0(n53[9]), 
          .S1(n53[10]));   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777_add_4_11.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1777_add_4_11.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1777_add_4_11.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1777_add_4_11.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1777_add_4_9 (.A0(pwm_freq_cntr[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n21864), .COUT(n21865), .S0(n53[7]), 
          .S1(n53[8]));   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777_add_4_9.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1777_add_4_9.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1777_add_4_9.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1777_add_4_9.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1777_add_4_7 (.A0(pwm_freq_cntr[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n21863), .COUT(n21864), .S0(n53[5]), 
          .S1(n53[6]));   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777_add_4_7.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1777_add_4_7.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1777_add_4_7.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1777_add_4_7.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1777_add_4_5 (.A0(pwm_freq_cntr[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n21862), .COUT(n21863), .S0(n53[3]), 
          .S1(n53[4]));   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777_add_4_5.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1777_add_4_5.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1777_add_4_5.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1777_add_4_5.INJECT1_1 = "NO";
    CCU2D equal_54_13_17466 (.A0(pwm_out_N_3154[3]), .B0(pwm_freq_cntr[3]), 
          .C0(pwm_out_N_3154[2]), .D0(pwm_freq_cntr[2]), .A1(pwm_out_N_3154[1]), 
          .B1(pwm_freq_cntr[1]), .C1(pwm_out_N_3154[0]), .D1(pwm_freq_cntr[0]), 
          .CIN(n21780), .COUT(n21781));
    defparam equal_54_13_17466.INIT0 = 16'h9009;
    defparam equal_54_13_17466.INIT1 = 16'h9009;
    defparam equal_54_13_17466.INJECT1_0 = "YES";
    defparam equal_54_13_17466.INJECT1_1 = "YES";
    CCU2D equal_52_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_out_N_3170[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n21774));   // c:/s_links/sources/pwm_controller.v(59[7:36])
    defparam equal_52_0.INIT0 = 16'hF000;
    defparam equal_52_0.INIT1 = 16'h5555;
    defparam equal_52_0.INJECT1_0 = "NO";
    defparam equal_52_0.INJECT1_1 = "YES";
    CCU2D pwm_freq_cntr_1777_add_4_3 (.A0(pwm_freq_cntr[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n21861), .COUT(n21862), .S0(n53[1]), 
          .S1(n53[2]));   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777_add_4_3.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1777_add_4_3.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1777_add_4_3.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1777_add_4_3.INJECT1_1 = "NO";
    CCU2D equal_54_11 (.A0(pwm_out_N_3154[7]), .B0(pwm_freq_cntr[7]), .C0(pwm_out_N_3154[6]), 
          .D0(pwm_freq_cntr[6]), .A1(pwm_out_N_3154[5]), .B1(pwm_freq_cntr[5]), 
          .C1(pwm_out_N_3154[4]), .D1(pwm_freq_cntr[4]), .CIN(n21779), 
          .COUT(n21780));
    defparam equal_54_11.INIT0 = 16'h9009;
    defparam equal_54_11.INIT1 = 16'h9009;
    defparam equal_54_11.INJECT1_0 = "YES";
    defparam equal_54_11.INJECT1_1 = "YES";
    CCU2D pwm_freq_cntr_1777_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_freq_cntr[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n21861), .S1(n53[0]));   // c:/s_links/sources/pwm_controller.v(71[22:42])
    defparam pwm_freq_cntr_1777_add_4_1.INIT0 = 16'hF000;
    defparam pwm_freq_cntr_1777_add_4_1.INIT1 = 16'h0555;
    defparam pwm_freq_cntr_1777_add_4_1.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1777_add_4_1.INJECT1_1 = "NO";
    CCU2D equal_54_9 (.A0(pwm_out_N_3154[11]), .B0(pwm_freq_cntr[11]), .C0(pwm_out_N_3154[10]), 
          .D0(pwm_freq_cntr[10]), .A1(pwm_out_N_3154[9]), .B1(pwm_freq_cntr[9]), 
          .C1(pwm_out_N_3154[8]), .D1(pwm_freq_cntr[8]), .CIN(n21778), 
          .COUT(n21779));
    defparam equal_54_9.INIT0 = 16'h9009;
    defparam equal_54_9.INIT1 = 16'h9009;
    defparam equal_54_9.INJECT1_0 = "YES";
    defparam equal_54_9.INJECT1_1 = "YES";
    CCU2D equal_54_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_out_N_3154[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n21778));   // c:/s_links/sources/pwm_controller.v(66[12:41])
    defparam equal_54_0.INIT0 = 16'hF000;
    defparam equal_54_0.INIT1 = 16'h5555;
    defparam equal_54_0.INJECT1_0 = "NO";
    defparam equal_54_0.INJECT1_1 = "YES";
    CCU2D sub_20_add_2_13 (.A0(pwm_freq[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n22032), .S0(pwm_out_N_3170[11]), .S1(pwm_out_N_3170[12]));   // c:/s_links/sources/pwm_controller.v(59[24:36])
    defparam sub_20_add_2_13.INIT0 = 16'h5555;
    defparam sub_20_add_2_13.INIT1 = 16'hffff;
    defparam sub_20_add_2_13.INJECT1_0 = "NO";
    defparam sub_20_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_20_add_2_11 (.A0(pwm_freq[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_freq[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22031), .COUT(n22032), .S0(pwm_out_N_3170[9]), 
          .S1(pwm_out_N_3170[10]));   // c:/s_links/sources/pwm_controller.v(59[24:36])
    defparam sub_20_add_2_11.INIT0 = 16'h5555;
    defparam sub_20_add_2_11.INIT1 = 16'h5555;
    defparam sub_20_add_2_11.INJECT1_0 = "NO";
    defparam sub_20_add_2_11.INJECT1_1 = "NO";
    CCU2D equal_52_13 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21777), 
          .S0(pwm_out_N_3169));
    defparam equal_52_13.INIT0 = 16'hFFFF;
    defparam equal_52_13.INIT1 = 16'h0000;
    defparam equal_52_13.INJECT1_0 = "NO";
    defparam equal_52_13.INJECT1_1 = "NO";
    CCU2D sub_20_add_2_9 (.A0(pwm_freq[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_freq[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22030), .COUT(n22031), .S0(pwm_out_N_3170[7]), 
          .S1(pwm_out_N_3170[8]));   // c:/s_links/sources/pwm_controller.v(59[24:36])
    defparam sub_20_add_2_9.INIT0 = 16'h5555;
    defparam sub_20_add_2_9.INIT1 = 16'h5555;
    defparam sub_20_add_2_9.INJECT1_0 = "NO";
    defparam sub_20_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_20_add_2_7 (.A0(pwm_freq[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_freq[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22029), .COUT(n22030), .S0(pwm_out_N_3170[5]), 
          .S1(pwm_out_N_3170[6]));   // c:/s_links/sources/pwm_controller.v(59[24:36])
    defparam sub_20_add_2_7.INIT0 = 16'h5555;
    defparam sub_20_add_2_7.INIT1 = 16'h5555;
    defparam sub_20_add_2_7.INJECT1_0 = "NO";
    defparam sub_20_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_20_add_2_5 (.A0(pwm_freq[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_freq[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22028), .COUT(n22029), .S0(pwm_out_N_3170[3]), 
          .S1(pwm_out_N_3170[4]));   // c:/s_links/sources/pwm_controller.v(59[24:36])
    defparam sub_20_add_2_5.INIT0 = 16'h5555;
    defparam sub_20_add_2_5.INIT1 = 16'h5555;
    defparam sub_20_add_2_5.INJECT1_0 = "NO";
    defparam sub_20_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_20_add_2_3 (.A0(pwm_freq[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_freq[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22027), .COUT(n22028), .S0(pwm_out_N_3170[1]), 
          .S1(pwm_out_N_3170[2]));   // c:/s_links/sources/pwm_controller.v(59[24:36])
    defparam sub_20_add_2_3.INIT0 = 16'h5555;
    defparam sub_20_add_2_3.INIT1 = 16'h5555;
    defparam sub_20_add_2_3.INJECT1_0 = "NO";
    defparam sub_20_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_20_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_freq[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n22027), .S1(pwm_out_N_3170[0]));   // c:/s_links/sources/pwm_controller.v(59[24:36])
    defparam sub_20_add_2_1.INIT0 = 16'hF000;
    defparam sub_20_add_2_1.INIT1 = 16'h5555;
    defparam sub_20_add_2_1.INJECT1_0 = "NO";
    defparam sub_20_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_24_add_2_13 (.A0(pwm_duty[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n22025), .S0(pwm_out_N_3154[11]), .S1(pwm_out_N_3154[12]));   // c:/s_links/sources/pwm_controller.v(66[29:41])
    defparam sub_24_add_2_13.INIT0 = 16'h5555;
    defparam sub_24_add_2_13.INIT1 = 16'hffff;
    defparam sub_24_add_2_13.INJECT1_0 = "NO";
    defparam sub_24_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_24_add_2_11 (.A0(pwm_duty[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22024), .COUT(n22025), .S0(pwm_out_N_3154[9]), 
          .S1(pwm_out_N_3154[10]));   // c:/s_links/sources/pwm_controller.v(66[29:41])
    defparam sub_24_add_2_11.INIT0 = 16'h5555;
    defparam sub_24_add_2_11.INIT1 = 16'h5555;
    defparam sub_24_add_2_11.INJECT1_0 = "NO";
    defparam sub_24_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_24_add_2_9 (.A0(pwm_duty[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22023), .COUT(n22024), .S0(pwm_out_N_3154[7]), 
          .S1(pwm_out_N_3154[8]));   // c:/s_links/sources/pwm_controller.v(66[29:41])
    defparam sub_24_add_2_9.INIT0 = 16'h5555;
    defparam sub_24_add_2_9.INIT1 = 16'h5555;
    defparam sub_24_add_2_9.INJECT1_0 = "NO";
    defparam sub_24_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_24_add_2_7 (.A0(pwm_duty[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22022), .COUT(n22023), .S0(pwm_out_N_3154[5]), 
          .S1(pwm_out_N_3154[6]));   // c:/s_links/sources/pwm_controller.v(66[29:41])
    defparam sub_24_add_2_7.INIT0 = 16'h5555;
    defparam sub_24_add_2_7.INIT1 = 16'h5555;
    defparam sub_24_add_2_7.INJECT1_0 = "NO";
    defparam sub_24_add_2_7.INJECT1_1 = "NO";
    CCU2D equal_52_13_17465 (.A0(pwm_out_N_3170[3]), .B0(pwm_freq_cntr[3]), 
          .C0(pwm_out_N_3170[2]), .D0(pwm_freq_cntr[2]), .A1(pwm_out_N_3170[1]), 
          .B1(pwm_freq_cntr[1]), .C1(pwm_out_N_3170[0]), .D1(pwm_freq_cntr[0]), 
          .CIN(n21776), .COUT(n21777));
    defparam equal_52_13_17465.INIT0 = 16'h9009;
    defparam equal_52_13_17465.INIT1 = 16'h9009;
    defparam equal_52_13_17465.INJECT1_0 = "YES";
    defparam equal_52_13_17465.INJECT1_1 = "YES";
    CCU2D sub_24_add_2_5 (.A0(pwm_duty[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22021), .COUT(n22022), .S0(pwm_out_N_3154[3]), 
          .S1(pwm_out_N_3154[4]));   // c:/s_links/sources/pwm_controller.v(66[29:41])
    defparam sub_24_add_2_5.INIT0 = 16'h5555;
    defparam sub_24_add_2_5.INIT1 = 16'h5555;
    defparam sub_24_add_2_5.INJECT1_0 = "NO";
    defparam sub_24_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_24_add_2_3 (.A0(pwm_duty[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22020), .COUT(n22021), .S0(pwm_out_N_3154[1]), 
          .S1(pwm_out_N_3154[2]));   // c:/s_links/sources/pwm_controller.v(66[29:41])
    defparam sub_24_add_2_3.INIT0 = 16'h5555;
    defparam sub_24_add_2_3.INIT1 = 16'h5555;
    defparam sub_24_add_2_3.INJECT1_0 = "NO";
    defparam sub_24_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_24_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_duty[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n22020), .S1(pwm_out_N_3154[0]));   // c:/s_links/sources/pwm_controller.v(66[29:41])
    defparam sub_24_add_2_1.INIT0 = 16'hF000;
    defparam sub_24_add_2_1.INIT1 = 16'h5555;
    defparam sub_24_add_2_1.INJECT1_0 = "NO";
    defparam sub_24_add_2_1.INJECT1_1 = "NO";
    CCU2D equal_52_11 (.A0(pwm_out_N_3170[7]), .B0(pwm_freq_cntr[7]), .C0(pwm_out_N_3170[6]), 
          .D0(pwm_freq_cntr[6]), .A1(pwm_out_N_3170[5]), .B1(pwm_freq_cntr[5]), 
          .C1(pwm_out_N_3170[4]), .D1(pwm_freq_cntr[4]), .CIN(n21775), 
          .COUT(n21776));
    defparam equal_52_11.INIT0 = 16'h9009;
    defparam equal_52_11.INIT1 = 16'h9009;
    defparam equal_52_11.INJECT1_0 = "YES";
    defparam equal_52_11.INJECT1_1 = "YES";
    CCU2D equal_52_9 (.A0(pwm_out_N_3170[11]), .B0(pwm_freq_cntr[11]), .C0(pwm_out_N_3170[10]), 
          .D0(pwm_freq_cntr[10]), .A1(pwm_out_N_3170[9]), .B1(pwm_freq_cntr[9]), 
          .C1(pwm_out_N_3170[8]), .D1(pwm_freq_cntr[8]), .CIN(n21774), 
          .COUT(n21775));
    defparam equal_52_9.INIT0 = 16'h9009;
    defparam equal_52_9.INIT1 = 16'h9009;
    defparam equal_52_9.INJECT1_0 = "YES";
    defparam equal_52_9.INJECT1_1 = "YES";
    LUT4 i1_4_lut (.A(n28249), .B(pwm_out_N_3169), .C(resetn_c), .D(n28243), 
         .Z(n25197)) /* synthesis lut_function=(A (B (C))+!A (B (C (D)))) */ ;   // c:/s_links/sources/pwm_controller.v(53[8] 75[4])
    defparam i1_4_lut.init = 16'hc080;
    LUT4 i1_4_lut_adj_863 (.A(pwm_duty[9]), .B(n28245), .C(n28231), .D(pwm_duty[0]), 
         .Z(n28249)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/pwm_controller.v(61[8:23])
    defparam i1_4_lut_adj_863.init = 16'hfffe;
    LUT4 i1_4_lut_adj_864 (.A(pwm_duty[1]), .B(pwm_duty[10]), .C(pwm_duty[11]), 
         .D(pwm_duty[4]), .Z(n28243)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/pwm_controller.v(61[8:23])
    defparam i1_4_lut_adj_864.init = 16'hfffe;
    LUT4 i1_4_lut_adj_865 (.A(pwm_duty[7]), .B(pwm_duty[3]), .C(pwm_duty[6]), 
         .D(pwm_duty[8]), .Z(n28245)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/pwm_controller.v(61[8:23])
    defparam i1_4_lut_adj_865.init = 16'hfffe;
    LUT4 i1_2_lut (.A(pwm_duty[2]), .B(pwm_duty[5]), .Z(n28231)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/pwm_controller.v(61[8:23])
    defparam i1_2_lut.init = 16'heeee;
    
endmodule
//
// Verilog Description of module \quad_decoder(DEV_ID=4) 
//

module \quad_decoder(DEV_ID=4)  (quad_count, clk, n30185, \quad_a[4] , 
            \quad_b[4] , \spi_data_out_r_39__N_1874[0] , \spi_data_out_r_39__N_2023[0] , 
            quad_buffer, \pin_intrpt[14] , clk_enable_683, \spi_data_r[0] , 
            quad_homing, clk_enable_684, spi_data_out_r_39__N_1914, spi_data_out_r_39__N_2103, 
            quad_set_valid_N_2098, \spi_data_out_r_39__N_1874[31] , \spi_data_out_r_39__N_2023[31] , 
            \spi_data_out_r_39__N_1874[30] , \spi_data_out_r_39__N_2023[30] , 
            \spi_data_out_r_39__N_1874[29] , \spi_data_out_r_39__N_2023[29] , 
            \spi_data_out_r_39__N_1874[28] , \spi_data_out_r_39__N_2023[28] , 
            \spi_data_out_r_39__N_1874[27] , \spi_data_out_r_39__N_2023[27] , 
            \spi_data_out_r_39__N_1874[26] , \spi_data_out_r_39__N_2023[26] , 
            \spi_data_out_r_39__N_1874[25] , \spi_data_out_r_39__N_2023[25] , 
            \spi_data_out_r_39__N_1874[24] , \spi_data_out_r_39__N_2023[24] , 
            \spi_data_out_r_39__N_1874[23] , \spi_data_out_r_39__N_2023[23] , 
            \spi_data_out_r_39__N_1874[22] , \spi_data_out_r_39__N_2023[22] , 
            \spi_data_out_r_39__N_1874[21] , \spi_data_out_r_39__N_2023[21] , 
            \spi_data_out_r_39__N_1874[20] , \spi_data_out_r_39__N_2023[20] , 
            \spi_data_out_r_39__N_1874[19] , \spi_data_out_r_39__N_2023[19] , 
            \spi_data_out_r_39__N_1874[18] , \spi_data_out_r_39__N_2023[18] , 
            \spi_data_out_r_39__N_1874[17] , \spi_data_out_r_39__N_2023[17] , 
            \spi_data_out_r_39__N_1874[16] , \spi_data_out_r_39__N_2023[16] , 
            \spi_data_out_r_39__N_1874[15] , \spi_data_out_r_39__N_2023[15] , 
            \spi_data_out_r_39__N_1874[14] , \spi_data_out_r_39__N_2023[14] , 
            \spi_data_out_r_39__N_1874[13] , \spi_data_out_r_39__N_2023[13] , 
            \spi_data_out_r_39__N_1874[12] , \spi_data_out_r_39__N_2023[12] , 
            \spi_data_out_r_39__N_1874[11] , \spi_data_out_r_39__N_2023[11] , 
            \spi_data_out_r_39__N_1874[10] , \spi_data_out_r_39__N_2023[10] , 
            \spi_data_out_r_39__N_1874[9] , \spi_data_out_r_39__N_2023[9] , 
            \spi_data_out_r_39__N_1874[8] , \spi_data_out_r_39__N_2023[8] , 
            \spi_data_out_r_39__N_1874[7] , \spi_data_out_r_39__N_2023[7] , 
            \spi_data_out_r_39__N_1874[6] , \spi_data_out_r_39__N_2023[6] , 
            \spi_data_out_r_39__N_1874[5] , \spi_data_out_r_39__N_2023[5] , 
            \spi_data_out_r_39__N_1874[4] , \spi_data_out_r_39__N_2023[4] , 
            \spi_data_out_r_39__N_1874[3] , \spi_data_out_r_39__N_2023[3] , 
            \spi_data_out_r_39__N_1874[2] , \spi_data_out_r_39__N_2023[2] , 
            \spi_data_out_r_39__N_1874[1] , \spi_data_out_r_39__N_2023[1] , 
            n1, \spi_data_r[1] , \spi_data_r[2] , \spi_data_r[3] , \spi_data_r[4] , 
            \spi_data_r[5] , \spi_data_r[6] , \spi_data_r[7] , \spi_data_r[8] , 
            \spi_data_r[9] , \spi_data_r[10] , \spi_data_r[11] , \spi_data_r[12] , 
            \spi_data_r[13] , \spi_data_r[14] , \spi_data_r[15] , \spi_data_r[16] , 
            \spi_data_r[17] , \spi_data_r[18] , \spi_data_r[19] , \spi_data_r[20] , 
            \spi_data_r[21] , \spi_data_r[22] , \spi_data_r[23] , \spi_data_r[24] , 
            \spi_data_r[25] , \spi_data_r[26] , \spi_data_r[27] , \spi_data_r[28] , 
            \spi_data_r[29] , \spi_data_r[30] , \spi_data_r[31] , GND_net, 
            resetn_c) /* synthesis syn_module_defined=1 */ ;
    output [31:0]quad_count;
    input clk;
    input n30185;
    input \quad_a[4] ;
    input \quad_b[4] ;
    output \spi_data_out_r_39__N_1874[0] ;
    input \spi_data_out_r_39__N_2023[0] ;
    output [31:0]quad_buffer;
    input \pin_intrpt[14] ;
    input clk_enable_683;
    input \spi_data_r[0] ;
    output [1:0]quad_homing;
    input clk_enable_684;
    output spi_data_out_r_39__N_1914;
    input spi_data_out_r_39__N_2103;
    input quad_set_valid_N_2098;
    output \spi_data_out_r_39__N_1874[31] ;
    input \spi_data_out_r_39__N_2023[31] ;
    output \spi_data_out_r_39__N_1874[30] ;
    input \spi_data_out_r_39__N_2023[30] ;
    output \spi_data_out_r_39__N_1874[29] ;
    input \spi_data_out_r_39__N_2023[29] ;
    output \spi_data_out_r_39__N_1874[28] ;
    input \spi_data_out_r_39__N_2023[28] ;
    output \spi_data_out_r_39__N_1874[27] ;
    input \spi_data_out_r_39__N_2023[27] ;
    output \spi_data_out_r_39__N_1874[26] ;
    input \spi_data_out_r_39__N_2023[26] ;
    output \spi_data_out_r_39__N_1874[25] ;
    input \spi_data_out_r_39__N_2023[25] ;
    output \spi_data_out_r_39__N_1874[24] ;
    input \spi_data_out_r_39__N_2023[24] ;
    output \spi_data_out_r_39__N_1874[23] ;
    input \spi_data_out_r_39__N_2023[23] ;
    output \spi_data_out_r_39__N_1874[22] ;
    input \spi_data_out_r_39__N_2023[22] ;
    output \spi_data_out_r_39__N_1874[21] ;
    input \spi_data_out_r_39__N_2023[21] ;
    output \spi_data_out_r_39__N_1874[20] ;
    input \spi_data_out_r_39__N_2023[20] ;
    output \spi_data_out_r_39__N_1874[19] ;
    input \spi_data_out_r_39__N_2023[19] ;
    output \spi_data_out_r_39__N_1874[18] ;
    input \spi_data_out_r_39__N_2023[18] ;
    output \spi_data_out_r_39__N_1874[17] ;
    input \spi_data_out_r_39__N_2023[17] ;
    output \spi_data_out_r_39__N_1874[16] ;
    input \spi_data_out_r_39__N_2023[16] ;
    output \spi_data_out_r_39__N_1874[15] ;
    input \spi_data_out_r_39__N_2023[15] ;
    output \spi_data_out_r_39__N_1874[14] ;
    input \spi_data_out_r_39__N_2023[14] ;
    output \spi_data_out_r_39__N_1874[13] ;
    input \spi_data_out_r_39__N_2023[13] ;
    output \spi_data_out_r_39__N_1874[12] ;
    input \spi_data_out_r_39__N_2023[12] ;
    output \spi_data_out_r_39__N_1874[11] ;
    input \spi_data_out_r_39__N_2023[11] ;
    output \spi_data_out_r_39__N_1874[10] ;
    input \spi_data_out_r_39__N_2023[10] ;
    output \spi_data_out_r_39__N_1874[9] ;
    input \spi_data_out_r_39__N_2023[9] ;
    output \spi_data_out_r_39__N_1874[8] ;
    input \spi_data_out_r_39__N_2023[8] ;
    output \spi_data_out_r_39__N_1874[7] ;
    input \spi_data_out_r_39__N_2023[7] ;
    output \spi_data_out_r_39__N_1874[6] ;
    input \spi_data_out_r_39__N_2023[6] ;
    output \spi_data_out_r_39__N_1874[5] ;
    input \spi_data_out_r_39__N_2023[5] ;
    output \spi_data_out_r_39__N_1874[4] ;
    input \spi_data_out_r_39__N_2023[4] ;
    output \spi_data_out_r_39__N_1874[3] ;
    input \spi_data_out_r_39__N_2023[3] ;
    output \spi_data_out_r_39__N_1874[2] ;
    input \spi_data_out_r_39__N_2023[2] ;
    output \spi_data_out_r_39__N_1874[1] ;
    input \spi_data_out_r_39__N_2023[1] ;
    input n1;
    input \spi_data_r[1] ;
    input \spi_data_r[2] ;
    input \spi_data_r[3] ;
    input \spi_data_r[4] ;
    input \spi_data_r[5] ;
    input \spi_data_r[6] ;
    input \spi_data_r[7] ;
    input \spi_data_r[8] ;
    input \spi_data_r[9] ;
    input \spi_data_r[10] ;
    input \spi_data_r[11] ;
    input \spi_data_r[12] ;
    input \spi_data_r[13] ;
    input \spi_data_r[14] ;
    input \spi_data_r[15] ;
    input \spi_data_r[16] ;
    input \spi_data_r[17] ;
    input \spi_data_r[18] ;
    input \spi_data_r[19] ;
    input \spi_data_r[20] ;
    input \spi_data_r[21] ;
    input \spi_data_r[22] ;
    input \spi_data_r[23] ;
    input \spi_data_r[24] ;
    input \spi_data_r[25] ;
    input \spi_data_r[26] ;
    input \spi_data_r[27] ;
    input \spi_data_r[28] ;
    input \spi_data_r[29] ;
    input \spi_data_r[30] ;
    input \spi_data_r[31] ;
    input GND_net;
    input resetn_c;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire \pin_intrpt[14]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[14] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    
    wire clk_enable_420, n8544;
    wire [2:0]quad_a_delayed;   // c:/s_links/sources/quad_decoder.v(34[20:34])
    wire [2:0]quad_b_delayed;   // c:/s_links/sources/quad_decoder.v(35[19:33])
    wire [31:0]quad_set;   // c:/s_links/sources/quad_decoder.v(39[31:39])
    
    wire quad_set_valid, n9697, n9695, n9693, n9691, n9689, n9687, 
        n9685, n9683, n9681, n9679, n9677, n9675, n9673, n9671, 
        n9669, n9667, n9665, n9663, n9661, n9659, n9657, n9655, 
        n9653, n9651, n9649, n9647, n9645, n9643, n9641, n9639, 
        n9637, n6, count_dir;
    wire [31:0]n3963;
    
    wire n5711, n22079, n22078, n22077, n22076, n22075, n22074, 
        n22073, n22072, n22071, n22070, n22069, n22068, n22067, 
        n22066, n22065, n22064;
    
    FD1P3AX quad_count_i0_i0 (.D(n8544), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i0.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i0 (.D(\quad_a[4] ), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i0.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i0 (.D(\quad_b[4] ), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_2023[0] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX quad_buffer_i0 (.D(quad_count[0]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i0.GSR = "DISABLED";
    FD1P3IX quad_set__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i0.GSR = "DISABLED";
    FD1P3IX quad_homing__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_684), .CD(n30185), 
            .CK(clk), .Q(quad_homing[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(62[8] 69[4])
    defparam quad_homing__i0.GSR = "DISABLED";
    FD1S3IX i39_391 (.D(spi_data_out_r_39__N_2103), .CK(clk), .CD(n30185), 
            .Q(spi_data_out_r_39__N_1914)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam i39_391.GSR = "DISABLED";
    FD1S3IX quad_set_valid_388 (.D(quad_set_valid_N_2098), .CK(clk), .CD(n30185), 
            .Q(quad_set_valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set_valid_388.GSR = "DISABLED";
    FD1S3AX quad_buffer_i31 (.D(quad_count[31]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i31.GSR = "DISABLED";
    FD1S3AX quad_buffer_i30 (.D(quad_count[30]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i30.GSR = "DISABLED";
    FD1S3AX quad_buffer_i29 (.D(quad_count[29]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i29.GSR = "DISABLED";
    FD1S3AX quad_buffer_i28 (.D(quad_count[28]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i28.GSR = "DISABLED";
    FD1S3AX quad_buffer_i27 (.D(quad_count[27]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i27.GSR = "DISABLED";
    FD1S3AX quad_buffer_i26 (.D(quad_count[26]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i26.GSR = "DISABLED";
    FD1S3AX quad_buffer_i25 (.D(quad_count[25]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i25.GSR = "DISABLED";
    FD1S3AX quad_buffer_i24 (.D(quad_count[24]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i24.GSR = "DISABLED";
    FD1S3AX quad_buffer_i23 (.D(quad_count[23]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i23.GSR = "DISABLED";
    FD1S3AX quad_buffer_i22 (.D(quad_count[22]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i22.GSR = "DISABLED";
    FD1S3AX quad_buffer_i21 (.D(quad_count[21]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i21.GSR = "DISABLED";
    FD1S3AX quad_buffer_i20 (.D(quad_count[20]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i20.GSR = "DISABLED";
    FD1S3AX quad_buffer_i19 (.D(quad_count[19]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i19.GSR = "DISABLED";
    FD1S3AX quad_buffer_i18 (.D(quad_count[18]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i18.GSR = "DISABLED";
    FD1S3AX quad_buffer_i17 (.D(quad_count[17]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i17.GSR = "DISABLED";
    FD1S3AX quad_buffer_i16 (.D(quad_count[16]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i16.GSR = "DISABLED";
    FD1S3AX quad_buffer_i15 (.D(quad_count[15]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i15.GSR = "DISABLED";
    FD1S3AX quad_buffer_i14 (.D(quad_count[14]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i14.GSR = "DISABLED";
    FD1S3AX quad_buffer_i13 (.D(quad_count[13]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i13.GSR = "DISABLED";
    FD1S3AX quad_buffer_i12 (.D(quad_count[12]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i12.GSR = "DISABLED";
    FD1S3AX quad_buffer_i11 (.D(quad_count[11]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i11.GSR = "DISABLED";
    FD1S3AX quad_buffer_i10 (.D(quad_count[10]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i10.GSR = "DISABLED";
    FD1S3AX quad_buffer_i9 (.D(quad_count[9]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i9.GSR = "DISABLED";
    FD1S3AX quad_buffer_i8 (.D(quad_count[8]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i8.GSR = "DISABLED";
    FD1S3AX quad_buffer_i7 (.D(quad_count[7]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i7.GSR = "DISABLED";
    FD1S3AX quad_buffer_i6 (.D(quad_count[6]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i6.GSR = "DISABLED";
    FD1S3AX quad_buffer_i5 (.D(quad_count[5]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i5.GSR = "DISABLED";
    FD1S3AX quad_buffer_i4 (.D(quad_count[4]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i4.GSR = "DISABLED";
    FD1S3AX quad_buffer_i3 (.D(quad_count[3]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i3.GSR = "DISABLED";
    FD1S3AX quad_buffer_i2 (.D(quad_count[2]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i2.GSR = "DISABLED";
    FD1S3AX quad_buffer_i1 (.D(quad_count[1]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_2023[31] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i31 (.D(\spi_data_out_r_39__N_2023[30] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i30 (.D(\spi_data_out_r_39__N_2023[29] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i29 (.D(\spi_data_out_r_39__N_2023[28] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i28 (.D(\spi_data_out_r_39__N_2023[27] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i27 (.D(\spi_data_out_r_39__N_2023[26] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i26 (.D(\spi_data_out_r_39__N_2023[25] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i25 (.D(\spi_data_out_r_39__N_2023[24] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i24 (.D(\spi_data_out_r_39__N_2023[23] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i23 (.D(\spi_data_out_r_39__N_2023[22] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i22 (.D(\spi_data_out_r_39__N_2023[21] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i21 (.D(\spi_data_out_r_39__N_2023[20] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i20 (.D(\spi_data_out_r_39__N_2023[19] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i19 (.D(\spi_data_out_r_39__N_2023[18] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i18 (.D(\spi_data_out_r_39__N_2023[17] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i17 (.D(\spi_data_out_r_39__N_2023[16] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i16 (.D(\spi_data_out_r_39__N_2023[15] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_2023[14] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_2023[13] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_2023[12] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_2023[11] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_2023[10] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_2023[9] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_2023[8] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_2023[7] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_2023[6] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_2023[5] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_2023[4] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_2023[3] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_2023[2] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_2023[1] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1874[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i2 (.D(quad_b_delayed[1]), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i2.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i1 (.D(quad_b_delayed[0]), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i1.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i2 (.D(quad_a_delayed[1]), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i2.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i1 (.D(quad_a_delayed[0]), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i1.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i31 (.D(n9697), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i31.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i30 (.D(n9695), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i30.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i29 (.D(n9693), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i29.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i28 (.D(n9691), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i28.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i27 (.D(n9689), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i27.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i26 (.D(n9687), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i26.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i25 (.D(n9685), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i25.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i24 (.D(n9683), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i24.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i23 (.D(n9681), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i23.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i22 (.D(n9679), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i22.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i21 (.D(n9677), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i21.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i20 (.D(n9675), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i20.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i19 (.D(n9673), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i19.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i18 (.D(n9671), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i18.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i17 (.D(n9669), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i17.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i16 (.D(n9667), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i16.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i15 (.D(n9665), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i15.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i14 (.D(n9663), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i14.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i13 (.D(n9661), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i13.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i12 (.D(n9659), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i12.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i11 (.D(n9657), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i11.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i10 (.D(n9655), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i10.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i9 (.D(n9653), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i9.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i8 (.D(n9651), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i8.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i7 (.D(n9649), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i7.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i6 (.D(n9647), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i6.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i5 (.D(n9645), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i5.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i4 (.D(n9643), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i4.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i3 (.D(n9641), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i3.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i2 (.D(n9639), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i1 (.D(n9637), .SP(clk_enable_420), .CK(clk), 
            .Q(quad_count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i1.GSR = "DISABLED";
    LUT4 i2_2_lut (.A(quad_b_delayed[1]), .B(quad_a_delayed[2]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(96[19:96])
    defparam i2_2_lut.init = 16'h6666;
    LUT4 i1_2_lut (.A(quad_a_delayed[1]), .B(quad_b_delayed[2]), .Z(count_dir)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(96[19:96])
    defparam i1_2_lut.init = 16'h6666;
    LUT4 i5373_4_lut (.A(n3963[31]), .B(quad_set[31]), .C(n5711), .D(n1), 
         .Z(n9697)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5373_4_lut.init = 16'hc0ca;
    FD1P3IX quad_set__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i1.GSR = "DISABLED";
    FD1P3IX quad_set__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i2.GSR = "DISABLED";
    FD1P3IX quad_set__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i3.GSR = "DISABLED";
    FD1P3IX quad_set__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i4.GSR = "DISABLED";
    FD1P3IX quad_set__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i5.GSR = "DISABLED";
    FD1P3IX quad_set__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i6.GSR = "DISABLED";
    FD1P3IX quad_set__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i7.GSR = "DISABLED";
    FD1P3IX quad_set__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i8.GSR = "DISABLED";
    FD1P3IX quad_set__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i9.GSR = "DISABLED";
    FD1P3IX quad_set__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i10.GSR = "DISABLED";
    FD1P3IX quad_set__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i11.GSR = "DISABLED";
    FD1P3IX quad_set__i12 (.D(\spi_data_r[12] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i12.GSR = "DISABLED";
    FD1P3IX quad_set__i13 (.D(\spi_data_r[13] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i13.GSR = "DISABLED";
    FD1P3IX quad_set__i14 (.D(\spi_data_r[14] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i14.GSR = "DISABLED";
    FD1P3IX quad_set__i15 (.D(\spi_data_r[15] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i15.GSR = "DISABLED";
    FD1P3IX quad_set__i16 (.D(\spi_data_r[16] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i16.GSR = "DISABLED";
    FD1P3IX quad_set__i17 (.D(\spi_data_r[17] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i17.GSR = "DISABLED";
    FD1P3IX quad_set__i18 (.D(\spi_data_r[18] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i18.GSR = "DISABLED";
    FD1P3IX quad_set__i19 (.D(\spi_data_r[19] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i19.GSR = "DISABLED";
    FD1P3IX quad_set__i20 (.D(\spi_data_r[20] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i20.GSR = "DISABLED";
    FD1P3IX quad_set__i21 (.D(\spi_data_r[21] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i21.GSR = "DISABLED";
    FD1P3IX quad_set__i22 (.D(\spi_data_r[22] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i22.GSR = "DISABLED";
    FD1P3IX quad_set__i23 (.D(\spi_data_r[23] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i23.GSR = "DISABLED";
    FD1P3IX quad_set__i24 (.D(\spi_data_r[24] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i24.GSR = "DISABLED";
    FD1P3IX quad_set__i25 (.D(\spi_data_r[25] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i25.GSR = "DISABLED";
    FD1P3IX quad_set__i26 (.D(\spi_data_r[26] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i26.GSR = "DISABLED";
    FD1P3IX quad_set__i27 (.D(\spi_data_r[27] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i27.GSR = "DISABLED";
    FD1P3IX quad_set__i28 (.D(\spi_data_r[28] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i28.GSR = "DISABLED";
    FD1P3IX quad_set__i29 (.D(\spi_data_r[29] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i29.GSR = "DISABLED";
    FD1P3IX quad_set__i30 (.D(\spi_data_r[30] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i30.GSR = "DISABLED";
    FD1P3IX quad_set__i31 (.D(\spi_data_r[31] ), .SP(clk_enable_683), .CD(n30185), 
            .CK(clk), .Q(quad_set[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i31.GSR = "DISABLED";
    FD1P3IX quad_homing__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_684), .CD(n30185), 
            .CK(clk), .Q(quad_homing[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(62[8] 69[4])
    defparam quad_homing__i1.GSR = "DISABLED";
    LUT4 i5371_4_lut (.A(n3963[30]), .B(quad_set[30]), .C(n5711), .D(n1), 
         .Z(n9695)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5371_4_lut.init = 16'hc0ca;
    CCU2D add_1369_33 (.A0(quad_count[30]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[31]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22079), .S0(n3963[30]), .S1(n3963[31]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_33.INIT0 = 16'h5569;
    defparam add_1369_33.INIT1 = 16'h5569;
    defparam add_1369_33.INJECT1_0 = "NO";
    defparam add_1369_33.INJECT1_1 = "NO";
    CCU2D add_1369_31 (.A0(quad_count[28]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[29]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22078), .COUT(n22079), .S0(n3963[28]), .S1(n3963[29]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_31.INIT0 = 16'h5569;
    defparam add_1369_31.INIT1 = 16'h5569;
    defparam add_1369_31.INJECT1_0 = "NO";
    defparam add_1369_31.INJECT1_1 = "NO";
    CCU2D add_1369_29 (.A0(quad_count[26]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[27]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22077), .COUT(n22078), .S0(n3963[26]), .S1(n3963[27]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_29.INIT0 = 16'h5569;
    defparam add_1369_29.INIT1 = 16'h5569;
    defparam add_1369_29.INJECT1_0 = "NO";
    defparam add_1369_29.INJECT1_1 = "NO";
    CCU2D add_1369_27 (.A0(quad_count[24]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[25]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22076), .COUT(n22077), .S0(n3963[24]), .S1(n3963[25]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_27.INIT0 = 16'h5569;
    defparam add_1369_27.INIT1 = 16'h5569;
    defparam add_1369_27.INJECT1_0 = "NO";
    defparam add_1369_27.INJECT1_1 = "NO";
    CCU2D add_1369_25 (.A0(quad_count[22]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[23]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22075), .COUT(n22076), .S0(n3963[22]), .S1(n3963[23]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_25.INIT0 = 16'h5569;
    defparam add_1369_25.INIT1 = 16'h5569;
    defparam add_1369_25.INJECT1_0 = "NO";
    defparam add_1369_25.INJECT1_1 = "NO";
    CCU2D add_1369_23 (.A0(quad_count[20]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[21]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22074), .COUT(n22075), .S0(n3963[20]), .S1(n3963[21]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_23.INIT0 = 16'h5569;
    defparam add_1369_23.INIT1 = 16'h5569;
    defparam add_1369_23.INJECT1_0 = "NO";
    defparam add_1369_23.INJECT1_1 = "NO";
    CCU2D add_1369_21 (.A0(quad_count[18]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[19]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22073), .COUT(n22074), .S0(n3963[18]), .S1(n3963[19]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_21.INIT0 = 16'h5569;
    defparam add_1369_21.INIT1 = 16'h5569;
    defparam add_1369_21.INJECT1_0 = "NO";
    defparam add_1369_21.INJECT1_1 = "NO";
    CCU2D add_1369_19 (.A0(quad_count[16]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[17]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22072), .COUT(n22073), .S0(n3963[16]), .S1(n3963[17]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_19.INIT0 = 16'h5569;
    defparam add_1369_19.INIT1 = 16'h5569;
    defparam add_1369_19.INJECT1_0 = "NO";
    defparam add_1369_19.INJECT1_1 = "NO";
    CCU2D add_1369_17 (.A0(quad_count[14]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[15]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22071), .COUT(n22072), .S0(n3963[14]), .S1(n3963[15]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_17.INIT0 = 16'h5569;
    defparam add_1369_17.INIT1 = 16'h5569;
    defparam add_1369_17.INJECT1_0 = "NO";
    defparam add_1369_17.INJECT1_1 = "NO";
    CCU2D add_1369_15 (.A0(quad_count[12]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[13]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22070), .COUT(n22071), .S0(n3963[12]), .S1(n3963[13]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_15.INIT0 = 16'h5569;
    defparam add_1369_15.INIT1 = 16'h5569;
    defparam add_1369_15.INJECT1_0 = "NO";
    defparam add_1369_15.INJECT1_1 = "NO";
    CCU2D add_1369_13 (.A0(quad_count[10]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[11]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22069), .COUT(n22070), .S0(n3963[10]), .S1(n3963[11]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_13.INIT0 = 16'h5569;
    defparam add_1369_13.INIT1 = 16'h5569;
    defparam add_1369_13.INJECT1_0 = "NO";
    defparam add_1369_13.INJECT1_1 = "NO";
    CCU2D add_1369_11 (.A0(quad_count[8]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[9]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22068), .COUT(n22069), .S0(n3963[8]), .S1(n3963[9]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_11.INIT0 = 16'h5569;
    defparam add_1369_11.INIT1 = 16'h5569;
    defparam add_1369_11.INJECT1_0 = "NO";
    defparam add_1369_11.INJECT1_1 = "NO";
    CCU2D add_1369_9 (.A0(quad_count[6]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[7]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22067), .COUT(n22068), .S0(n3963[6]), .S1(n3963[7]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_9.INIT0 = 16'h5569;
    defparam add_1369_9.INIT1 = 16'h5569;
    defparam add_1369_9.INJECT1_0 = "NO";
    defparam add_1369_9.INJECT1_1 = "NO";
    CCU2D add_1369_7 (.A0(quad_count[4]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[5]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22066), .COUT(n22067), .S0(n3963[4]), .S1(n3963[5]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_7.INIT0 = 16'h5569;
    defparam add_1369_7.INIT1 = 16'h5569;
    defparam add_1369_7.INJECT1_0 = "NO";
    defparam add_1369_7.INJECT1_1 = "NO";
    CCU2D add_1369_5 (.A0(quad_count[2]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[3]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22065), .COUT(n22066), .S0(n3963[2]), .S1(n3963[3]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_5.INIT0 = 16'h5569;
    defparam add_1369_5.INIT1 = 16'h5569;
    defparam add_1369_5.INJECT1_0 = "NO";
    defparam add_1369_5.INJECT1_1 = "NO";
    CCU2D add_1369_3 (.A0(quad_count[0]), .B0(count_dir), .C0(n6), .D0(count_dir), 
          .A1(quad_count[1]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22064), .COUT(n22065), .S0(n3963[0]), .S1(n3963[1]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_3.INIT0 = 16'h5665;
    defparam add_1369_3.INIT1 = 16'h5569;
    defparam add_1369_3.INJECT1_0 = "NO";
    defparam add_1369_3.INJECT1_1 = "NO";
    CCU2D add_1369_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quad_a_delayed[2]), .B1(quad_b_delayed[1]), .C1(quad_b_delayed[2]), 
          .D1(quad_a_delayed[1]), .COUT(n22064));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1369_1.INIT0 = 16'hF000;
    defparam add_1369_1.INIT1 = 16'h0990;
    defparam add_1369_1.INJECT1_0 = "NO";
    defparam add_1369_1.INJECT1_1 = "NO";
    LUT4 i24190_2_lut (.A(resetn_c), .B(quad_homing[1]), .Z(clk_enable_420)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i24190_2_lut.init = 16'h7777;
    LUT4 i4220_4_lut (.A(n3963[0]), .B(quad_set[0]), .C(n5711), .D(n1), 
         .Z(n8544)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4220_4_lut.init = 16'hc0ca;
    LUT4 i1_4_lut (.A(quad_homing[0]), .B(quad_homing[1]), .C(quad_set_valid), 
         .D(resetn_c), .Z(n5711)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut.init = 16'h1000;
    LUT4 i5369_4_lut (.A(n3963[29]), .B(quad_set[29]), .C(n5711), .D(n1), 
         .Z(n9693)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5369_4_lut.init = 16'hc0ca;
    LUT4 i5367_4_lut (.A(n3963[28]), .B(quad_set[28]), .C(n5711), .D(n1), 
         .Z(n9691)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5367_4_lut.init = 16'hc0ca;
    LUT4 i5365_4_lut (.A(n3963[27]), .B(quad_set[27]), .C(n5711), .D(n1), 
         .Z(n9689)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5365_4_lut.init = 16'hc0ca;
    LUT4 i5363_4_lut (.A(n3963[26]), .B(quad_set[26]), .C(n5711), .D(n1), 
         .Z(n9687)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5363_4_lut.init = 16'hc0ca;
    LUT4 i5361_4_lut (.A(n3963[25]), .B(quad_set[25]), .C(n5711), .D(n1), 
         .Z(n9685)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5361_4_lut.init = 16'hc0ca;
    LUT4 i5359_4_lut (.A(n3963[24]), .B(quad_set[24]), .C(n5711), .D(n1), 
         .Z(n9683)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5359_4_lut.init = 16'hc0ca;
    LUT4 i5357_4_lut (.A(n3963[23]), .B(quad_set[23]), .C(n5711), .D(n1), 
         .Z(n9681)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5357_4_lut.init = 16'hc0ca;
    LUT4 i5355_4_lut (.A(n3963[22]), .B(quad_set[22]), .C(n5711), .D(n1), 
         .Z(n9679)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5355_4_lut.init = 16'hc0ca;
    LUT4 i5353_4_lut (.A(n3963[21]), .B(quad_set[21]), .C(n5711), .D(n1), 
         .Z(n9677)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5353_4_lut.init = 16'hc0ca;
    LUT4 i5351_4_lut (.A(n3963[20]), .B(quad_set[20]), .C(n5711), .D(n1), 
         .Z(n9675)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5351_4_lut.init = 16'hc0ca;
    LUT4 i5349_4_lut (.A(n3963[19]), .B(quad_set[19]), .C(n5711), .D(n1), 
         .Z(n9673)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5349_4_lut.init = 16'hc0ca;
    LUT4 i5347_4_lut (.A(n3963[18]), .B(quad_set[18]), .C(n5711), .D(n1), 
         .Z(n9671)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5347_4_lut.init = 16'hc0ca;
    LUT4 i5345_4_lut (.A(n3963[17]), .B(quad_set[17]), .C(n5711), .D(n1), 
         .Z(n9669)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5345_4_lut.init = 16'hc0ca;
    LUT4 i5343_4_lut (.A(n3963[16]), .B(quad_set[16]), .C(n5711), .D(n1), 
         .Z(n9667)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5343_4_lut.init = 16'hc0ca;
    LUT4 i5341_4_lut (.A(n3963[15]), .B(quad_set[15]), .C(n5711), .D(n1), 
         .Z(n9665)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5341_4_lut.init = 16'hc0ca;
    LUT4 i5339_4_lut (.A(n3963[14]), .B(quad_set[14]), .C(n5711), .D(n1), 
         .Z(n9663)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5339_4_lut.init = 16'hc0ca;
    LUT4 i5337_4_lut (.A(n3963[13]), .B(quad_set[13]), .C(n5711), .D(n1), 
         .Z(n9661)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5337_4_lut.init = 16'hc0ca;
    LUT4 i5335_4_lut (.A(n3963[12]), .B(quad_set[12]), .C(n5711), .D(n1), 
         .Z(n9659)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5335_4_lut.init = 16'hc0ca;
    LUT4 i5333_4_lut (.A(n3963[11]), .B(quad_set[11]), .C(n5711), .D(n1), 
         .Z(n9657)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5333_4_lut.init = 16'hc0ca;
    LUT4 i5331_4_lut (.A(n3963[10]), .B(quad_set[10]), .C(n5711), .D(n1), 
         .Z(n9655)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5331_4_lut.init = 16'hc0ca;
    LUT4 i5329_4_lut (.A(n3963[9]), .B(quad_set[9]), .C(n5711), .D(n1), 
         .Z(n9653)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5329_4_lut.init = 16'hc0ca;
    LUT4 i5327_4_lut (.A(n3963[8]), .B(quad_set[8]), .C(n5711), .D(n1), 
         .Z(n9651)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5327_4_lut.init = 16'hc0ca;
    LUT4 i5325_4_lut (.A(n3963[7]), .B(quad_set[7]), .C(n5711), .D(n1), 
         .Z(n9649)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5325_4_lut.init = 16'hc0ca;
    LUT4 i5323_4_lut (.A(n3963[6]), .B(quad_set[6]), .C(n5711), .D(n1), 
         .Z(n9647)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5323_4_lut.init = 16'hc0ca;
    LUT4 i5321_4_lut (.A(n3963[5]), .B(quad_set[5]), .C(n5711), .D(n1), 
         .Z(n9645)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5321_4_lut.init = 16'hc0ca;
    LUT4 i5319_4_lut (.A(n3963[4]), .B(quad_set[4]), .C(n5711), .D(n1), 
         .Z(n9643)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5319_4_lut.init = 16'hc0ca;
    LUT4 i5317_4_lut (.A(n3963[3]), .B(quad_set[3]), .C(n5711), .D(n1), 
         .Z(n9641)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5317_4_lut.init = 16'hc0ca;
    LUT4 i5315_4_lut (.A(n3963[2]), .B(quad_set[2]), .C(n5711), .D(n1), 
         .Z(n9639)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5315_4_lut.init = 16'hc0ca;
    LUT4 i5313_4_lut (.A(n3963[1]), .B(quad_set[1]), .C(n5711), .D(n1), 
         .Z(n9637)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5313_4_lut.init = 16'hc0ca;
    
endmodule
//
// Verilog Description of module \rs232(DEV_ID=4,UART_ADDRESS_WIDTH=4) 
//

module \rs232(DEV_ID=4,UART_ADDRESS_WIDTH=4)  (n28340, n24066, n28328, 
            quad_set_valid_N_2333, spi_addr_r, n30214, n25643, n30210, 
            mode, clk, clk_enable_253, n30185, \spi_data_r[0] , \spi_cmd_r[0] , 
            n26107, n26621, n26207, n30071, \spi_cmd_r[5] , n28476, 
            n26819, n30144, n26821, \spi_cmd_r[3] , n30155, n28260, 
            n30044, n25941, n18440, n30213, n25979, resetn_c, n30122, 
            \uart_slot_en[0] , \uart_slot_en[2] , \uart_slot_en[1] , TX_IN_N_6565, 
            n25739, UC_TXD0_c, n30180, n7164, n26633, n23916, n23526, 
            n30004, n26947, \spi_cmd_r[2] , n30199, n30031) /* synthesis syn_module_defined=1 */ ;
    output n28340;
    input n24066;
    input n28328;
    output quad_set_valid_N_2333;
    input [7:0]spi_addr_r;
    input n30214;
    input n25643;
    input n30210;
    output mode;
    input clk;
    input clk_enable_253;
    input n30185;
    input \spi_data_r[0] ;
    input \spi_cmd_r[0] ;
    input n26107;
    output n26621;
    output n26207;
    output n30071;
    input \spi_cmd_r[5] ;
    output n28476;
    input n26819;
    input n30144;
    output n26821;
    input \spi_cmd_r[3] ;
    output n30155;
    output n28260;
    input n30044;
    output n25941;
    input n18440;
    input n30213;
    output n25979;
    input resetn_c;
    input n30122;
    input \uart_slot_en[0] ;
    input \uart_slot_en[2] ;
    input \uart_slot_en[1] ;
    output TX_IN_N_6565;
    output n25739;
    input UC_TXD0_c;
    input n30180;
    output n7164;
    output n26633;
    input n23916;
    input n23526;
    output n30004;
    output n26947;
    input \spi_cmd_r[2] ;
    input n30199;
    output n30031;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    
    wire n25653, n28288, n28478, n25929, n25967, n25727, n28454, 
        n26943, n26931;
    
    LUT4 i1_4_lut (.A(n28340), .B(n24066), .C(n25653), .D(n28328), .Z(quad_set_valid_N_2333)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_adj_852 (.A(spi_addr_r[4]), .B(n30214), .C(n25643), 
         .D(n30210), .Z(n25653)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_852.init = 16'h1000;
    FD1P3IX mode_26 (.D(\spi_data_r[0] ), .SP(clk_enable_253), .CD(n30185), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=541, LSE_RLINE=561 */ ;   // c:/s_links/sources/rs232.v(39[8] 47[4])
    defparam mode_26.GSR = "DISABLED";
    LUT4 i23638_2_lut (.A(spi_addr_r[1]), .B(\spi_cmd_r[0] ), .Z(n28340)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23638_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_853 (.A(n26107), .B(n26621), .C(spi_addr_r[0]), 
         .D(n30214), .Z(n26207)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_853.init = 16'h0004;
    LUT4 i23754_2_lut_rep_671_3_lut (.A(spi_addr_r[5]), .B(spi_addr_r[7]), 
         .C(spi_addr_r[0]), .Z(n30071)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i23754_2_lut_rep_671_3_lut.init = 16'hfefe;
    LUT4 i23774_3_lut_4_lut (.A(spi_addr_r[5]), .B(spi_addr_r[7]), .C(\spi_cmd_r[5] ), 
         .D(spi_addr_r[6]), .Z(n28476)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23774_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_854 (.A(n26819), .B(n30144), .C(n28288), .D(spi_addr_r[3]), 
         .Z(n26821)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_854.init = 16'h0002;
    LUT4 i23586_2_lut (.A(\spi_cmd_r[3] ), .B(spi_addr_r[5]), .Z(n28288)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23586_2_lut.init = 16'heeee;
    LUT4 i23668_2_lut_rep_755 (.A(spi_addr_r[5]), .B(spi_addr_r[7]), .Z(n30155)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23668_2_lut_rep_755.init = 16'heeee;
    LUT4 i23559_2_lut (.A(spi_addr_r[1]), .B(spi_addr_r[7]), .Z(n28260)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23559_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_855 (.A(n28478), .B(n30044), .C(n30155), .D(n25929), 
         .Z(n25941)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_855.init = 16'h0400;
    LUT4 i1_4_lut_adj_856 (.A(n28478), .B(n18440), .C(n25967), .D(n30213), 
         .Z(n25979)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_856.init = 16'h0010;
    LUT4 i1_3_lut (.A(spi_addr_r[5]), .B(spi_addr_r[2]), .C(resetn_c), 
         .Z(n25967)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4040;
    LUT4 i3_4_lut (.A(n30122), .B(\uart_slot_en[0] ), .C(\uart_slot_en[2] ), 
         .D(\uart_slot_en[1] ), .Z(TX_IN_N_6565)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i3_4_lut.init = 16'h0020;
    LUT4 i1_4_lut_adj_857 (.A(n28478), .B(n30044), .C(n25727), .D(n30213), 
         .Z(n25739)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_adj_857.init = 16'h0040;
    LUT4 Select_2826_i3_3_lut (.A(UC_TXD0_c), .B(n30180), .C(TX_IN_N_6565), 
         .Z(n7164)) /* synthesis lut_function=(A ((C)+!B)+!A !(B)) */ ;
    defparam Select_2826_i3_3_lut.init = 16'hb3b3;
    LUT4 i1_4_lut_adj_858 (.A(n28454), .B(n18440), .C(n26621), .D(n30144), 
         .Z(n26633)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_858.init = 16'h0010;
    LUT4 i23752_3_lut (.A(spi_addr_r[3]), .B(spi_addr_r[0]), .C(spi_addr_r[5]), 
         .Z(n28454)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i23752_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut (.A(spi_addr_r[7]), .B(spi_addr_r[2]), .Z(n26621)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i1_3_lut_rep_604 (.A(n23916), .B(n23526), .C(n26207), .Z(n30004)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_rep_604.init = 16'h8080;
    LUT4 i1_2_lut_3_lut (.A(spi_addr_r[2]), .B(\spi_cmd_r[3] ), .C(spi_addr_r[4]), 
         .Z(n25929)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_3_lut_adj_859 (.A(spi_addr_r[2]), .B(\spi_cmd_r[3] ), 
         .C(spi_addr_r[5]), .Z(n25727)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_adj_859.init = 16'h0808;
    LUT4 i23776_3_lut (.A(spi_addr_r[3]), .B(spi_addr_r[0]), .C(spi_addr_r[6]), 
         .Z(n28478)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i23776_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_860 (.A(n26943), .B(n18440), .C(spi_addr_r[0]), 
         .D(n28260), .Z(n26947)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_860.init = 16'h0002;
    LUT4 i1_4_lut_adj_861 (.A(n30144), .B(spi_addr_r[3]), .C(n26931), 
         .D(\spi_cmd_r[0] ), .Z(n26943)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_861.init = 16'h0010;
    LUT4 i1_3_lut_adj_862 (.A(spi_addr_r[5]), .B(spi_addr_r[2]), .C(\spi_cmd_r[2] ), 
         .Z(n26931)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut_adj_862.init = 16'h4040;
    LUT4 i1_3_lut_rep_631 (.A(n26633), .B(n23916), .C(n30199), .Z(n30031)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_rep_631.init = 16'h8080;
    
endmodule
//
// Verilog Description of module \stepper(DEV_ID=2,UART_ADDRESS_WIDTH=4) 
//

module \stepper(DEV_ID=2,UART_ADDRESS_WIDTH=4)  (clk, clk_1MHz, n30185, 
            GND_net, pin_io_c_28, reset_r, clk_enable_23, n29996, 
            resetn_c, n30110, spi_data_out_r_39__N_4511, clk_enable_686, 
            \spi_data_r[0] , n47, spi_data_out_r_39__N_4551, spi_data_out_r_39__N_4848, 
            digital_output_r, clk_enable_259, n28556, \quad_homing[0] , 
            pin_io_c_24, n25881, \spi_data_r[1] , \mode[2] , \spi_data_r[2] , 
            NSL, n5, UC_TXD0_c, OW_ID_N_4804, n9, \uart_slot_en[0] , 
            \uart_slot_en[1] , pin_io_out_29, \quad_b[2] , \quad_a[2] , 
            pin_io_c_23, \pin_intrpt[7] , n30095, OW_ID_N_4810, pin_io_c_22, 
            \pin_intrpt[6] , \pin_intrpt[8] , n7273, ENC_O_N_4812) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input clk_1MHz;
    input n30185;
    input GND_net;
    input pin_io_c_28;
    output reset_r;
    input clk_enable_23;
    input n29996;
    input resetn_c;
    output n30110;
    output [39:0]spi_data_out_r_39__N_4511;
    input clk_enable_686;
    input \spi_data_r[0] ;
    input n47;
    output spi_data_out_r_39__N_4551;
    input spi_data_out_r_39__N_4848;
    output digital_output_r;
    input clk_enable_259;
    input n28556;
    input \quad_homing[0] ;
    input pin_io_c_24;
    output n25881;
    input \spi_data_r[1] ;
    output \mode[2] ;
    input \spi_data_r[2] ;
    output NSL;
    output n5;
    input UC_TXD0_c;
    output OW_ID_N_4804;
    input n9;
    input \uart_slot_en[0] ;
    input \uart_slot_en[1] ;
    input pin_io_out_29;
    output \quad_b[2] ;
    output \quad_a[2] ;
    input pin_io_c_23;
    output \pin_intrpt[7] ;
    output n30095;
    output OW_ID_N_4810;
    input pin_io_c_22;
    output \pin_intrpt[6] ;
    output \pin_intrpt[8] ;
    output n7273;
    output ENC_O_N_4812;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire clk_1MHz /* synthesis SET_AS_NETWORK=clk_1MHz, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(136[6:14])
    wire \pin_intrpt[8]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[8] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    wire [51:0]SLO;   // c:/s_links/sources/slot_cards/stepper.v(63[12:15])
    
    wire clk_enable_1135, n12391, MA_Temp, clk_1MHz_enable_1, MA_Temp_N_4830;
    wire [7:0]Cnt;   // c:/s_links/sources/slot_cards/stepper.v(62[11:14])
    
    wire n30202, n18578;
    wire [11:0]n93;
    wire [11:0]n53;
    
    wire prev_MA_Temp, n30100, n30099, n18664, clk_1MHz_enable_66, 
        prev_MA;
    wire [39:0]spi_data_out_r_39__N_4762;
    
    wire n18666, n28318, n30068, n28588;
    wire [2:0]mode;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    wire [51:0]SLO_buf;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire clk_1MHz_enable_64;
    wire [7:0]n199;
    
    wire SLO_buf_51__N_4701;
    wire [31:0]n153;
    wire [11:0]Cnt_NSL;   // c:/s_links/sources/slot_cards/stepper.v(61[12:19])
    
    wire n30040, n30003, NSL_N_4843, n28587, n30048, n26383, n4, 
        n21944, n21943, n21942, n21941, n21933, n21932, n21931, 
        n21930, n21929, n21928, n30097, OW_ID_N_4805, n28330, n30037, 
        n30215, n30152, n24971;
    
    FD1P3IX SLO__i25 (.D(SLO[23]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i25.GSR = "DISABLED";
    FD1P3IX MA_Temp_483 (.D(MA_Temp_N_4830), .SP(clk_1MHz_enable_1), .CD(n30185), 
            .CK(clk_1MHz), .Q(MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam MA_Temp_483.GSR = "DISABLED";
    FD1P3IX SLO__i26 (.D(SLO[24]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i26.GSR = "DISABLED";
    FD1P3IX SLO__i1 (.D(pin_io_c_28), .SP(clk_enable_1135), .CD(GND_net), 
            .CK(clk), .Q(SLO[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i1.GSR = "DISABLED";
    FD1P3IX SLO__i27 (.D(SLO[25]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i27.GSR = "DISABLED";
    FD1P3IX reset_r_491 (.D(n29996), .SP(clk_enable_23), .CD(n30185), 
            .CK(clk), .Q(reset_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam reset_r_491.GSR = "DISABLED";
    FD1P3IX SLO__i28 (.D(SLO[26]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i28.GSR = "DISABLED";
    FD1P3IX SLO__i29 (.D(SLO[27]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i29.GSR = "DISABLED";
    FD1P3IX SLO__i30 (.D(SLO[28]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i30.GSR = "DISABLED";
    FD1P3IX SLO__i2 (.D(SLO[0]), .SP(clk_enable_1135), .CD(GND_net), .CK(clk), 
            .Q(SLO[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i2.GSR = "DISABLED";
    FD1P3IX SLO__i3 (.D(SLO[1]), .SP(clk_enable_1135), .CD(GND_net), .CK(clk), 
            .Q(SLO[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i3.GSR = "DISABLED";
    FD1P3IX SLO__i4 (.D(SLO[2]), .SP(clk_enable_1135), .CD(GND_net), .CK(clk), 
            .Q(SLO[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i4.GSR = "DISABLED";
    FD1P3IX SLO__i31 (.D(SLO[29]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i31.GSR = "DISABLED";
    LUT4 i14251_2_lut_4_lut (.A(Cnt[0]), .B(n30202), .C(Cnt[1]), .D(Cnt[4]), 
         .Z(n18578)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(107[15:23])
    defparam i14251_2_lut_4_lut.init = 16'hec00;
    FD1P3IX SLO__i5 (.D(SLO[3]), .SP(clk_enable_1135), .CD(GND_net), .CK(clk), 
            .Q(SLO[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i5.GSR = "DISABLED";
    FD1P3IX SLO__i6 (.D(SLO[4]), .SP(clk_enable_1135), .CD(GND_net), .CK(clk), 
            .Q(SLO[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i6.GSR = "DISABLED";
    FD1P3IX SLO__i7 (.D(SLO[5]), .SP(clk_enable_1135), .CD(GND_net), .CK(clk), 
            .Q(SLO[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i7.GSR = "DISABLED";
    FD1P3IX SLO__i8 (.D(SLO[6]), .SP(clk_enable_1135), .CD(GND_net), .CK(clk), 
            .Q(SLO[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i8.GSR = "DISABLED";
    FD1P3IX SLO__i9 (.D(SLO[7]), .SP(clk_enable_1135), .CD(GND_net), .CK(clk), 
            .Q(SLO[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i9.GSR = "DISABLED";
    FD1P3IX SLO__i10 (.D(SLO[8]), .SP(clk_enable_1135), .CD(GND_net), 
            .CK(clk), .Q(SLO[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i10.GSR = "DISABLED";
    FD1P3IX SLO__i32 (.D(SLO[30]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i32.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1780__i0 (.D(n53[0]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780__i0.GSR = "DISABLED";
    FD1P3IX SLO__i33 (.D(SLO[31]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i33.GSR = "DISABLED";
    FD1P3IX SLO__i11 (.D(SLO[9]), .SP(clk_enable_1135), .CD(GND_net), 
            .CK(clk), .Q(SLO[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i11.GSR = "DISABLED";
    FD1P3IX SLO__i12 (.D(SLO[10]), .SP(clk_enable_1135), .CD(GND_net), 
            .CK(clk), .Q(SLO[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i12.GSR = "DISABLED";
    FD1P3IX SLO__i34 (.D(SLO[32]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i34.GSR = "DISABLED";
    FD1P3IX SLO__i13 (.D(SLO[11]), .SP(clk_enable_1135), .CD(GND_net), 
            .CK(clk), .Q(SLO[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i13.GSR = "DISABLED";
    FD1P3IX SLO__i14 (.D(SLO[12]), .SP(clk_enable_1135), .CD(GND_net), 
            .CK(clk), .Q(SLO[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i14.GSR = "DISABLED";
    FD1P3IX SLO__i15 (.D(SLO[13]), .SP(clk_enable_1135), .CD(GND_net), 
            .CK(clk), .Q(SLO[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i15.GSR = "DISABLED";
    FD1P3IX SLO__i16 (.D(SLO[14]), .SP(clk_enable_1135), .CD(GND_net), 
            .CK(clk), .Q(SLO[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i16.GSR = "DISABLED";
    FD1P3IX SLO__i35 (.D(SLO[33]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i35.GSR = "DISABLED";
    FD1P3IX SLO__i17 (.D(SLO[15]), .SP(clk_enable_1135), .CD(GND_net), 
            .CK(clk), .Q(SLO[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i17.GSR = "DISABLED";
    FD1P3IX SLO__i18 (.D(SLO[16]), .SP(clk_enable_1135), .CD(GND_net), 
            .CK(clk), .Q(SLO[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i18.GSR = "DISABLED";
    FD1S3AX prev_MA_Temp_487 (.D(MA_Temp), .CK(clk), .Q(prev_MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam prev_MA_Temp_487.GSR = "DISABLED";
    LUT4 i14052_3_lut_4_lut (.A(n30100), .B(n30099), .C(resetn_c), .D(n18664), 
         .Z(clk_1MHz_enable_66)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i14052_3_lut_4_lut.init = 16'h70f0;
    FD1S3AX prev_MA_489 (.D(n30110), .CK(clk), .Q(prev_MA)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam prev_MA_489.GSR = "DISABLED";
    FD1P3IX SLO__i36 (.D(SLO[34]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i36.GSR = "DISABLED";
    FD1P3IX SLO__i19 (.D(SLO[17]), .SP(clk_enable_1135), .CD(GND_net), 
            .CK(clk), .Q(SLO[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i19.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i0 (.D(spi_data_out_r_39__N_4762[0]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i0.GSR = "DISABLED";
    FD1P3IX SLO__i20 (.D(SLO[18]), .SP(clk_enable_1135), .CD(GND_net), 
            .CK(clk), .Q(SLO[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i20.GSR = "DISABLED";
    FD1P3IX SLO__i21 (.D(SLO[19]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i21.GSR = "DISABLED";
    FD1P3IX SLO__i22 (.D(SLO[20]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i22.GSR = "DISABLED";
    FD1P3IX SLO__i23 (.D(SLO[21]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i23.GSR = "DISABLED";
    FD1P3IX SLO__i37 (.D(SLO[35]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i37.GSR = "DISABLED";
    LUT4 i23895_1_lut_4_lut (.A(MA_Temp), .B(n18666), .C(n28318), .D(n30068), 
         .Z(n28588)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A (B+((D)+!C)))) */ ;
    defparam i23895_1_lut_4_lut.init = 16'h2212;
    FD1P3IX mode__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_686), .CD(n30185), 
            .CK(clk), .Q(mode[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i0.GSR = "DISABLED";
    FD1P3IX SLO__i38 (.D(SLO[36]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i38.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i39 (.D(SLO_buf[13]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i39.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i38 (.D(SLO_buf[12]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i38.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i37 (.D(SLO_buf[11]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i37.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i36 (.D(SLO_buf[10]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i36.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i35 (.D(spi_data_out_r_39__N_4762[35]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i35.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i34 (.D(spi_data_out_r_39__N_4762[34]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i34.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i33 (.D(spi_data_out_r_39__N_4762[33]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i33.GSR = "DISABLED";
    FD1P3IX SLO__i39 (.D(SLO[37]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i39.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(spi_data_out_r_39__N_4762[32]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i31 (.D(SLO_buf[45]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i30 (.D(SLO_buf[44]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i29 (.D(SLO_buf[43]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i28 (.D(SLO_buf[42]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i27 (.D(SLO_buf[41]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i26 (.D(SLO_buf[40]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i25 (.D(SLO_buf[39]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i24 (.D(SLO_buf[38]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i23 (.D(SLO_buf[37]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i22 (.D(SLO_buf[36]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i21 (.D(SLO_buf[35]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i20 (.D(SLO_buf[34]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i19 (.D(SLO_buf[33]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i18 (.D(SLO_buf[32]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i17 (.D(SLO_buf[31]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i16 (.D(SLO_buf[30]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4511[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1P3IX SLO__i40 (.D(SLO[38]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i40.GSR = "DISABLED";
    FD1P3IX Cnt__i0 (.D(n199[0]), .SP(clk_1MHz_enable_64), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i0.GSR = "DISABLED";
    FD1P3IX SLO__i41 (.D(SLO[39]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i41.GSR = "DISABLED";
    FD1P3IX SLO__i42 (.D(SLO[40]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i42.GSR = "DISABLED";
    FD1P3AX SLO_buf__i1 (.D(SLO[0]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(spi_data_out_r_39__N_4762[15]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(spi_data_out_r_39__N_4762[14]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(spi_data_out_r_39__N_4762[13]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(spi_data_out_r_39__N_4762[12]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(spi_data_out_r_39__N_4762[11]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(spi_data_out_r_39__N_4762[10]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(spi_data_out_r_39__N_4762[9]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(spi_data_out_r_39__N_4762[8]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(spi_data_out_r_39__N_4762[7]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(spi_data_out_r_39__N_4762[6]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(spi_data_out_r_39__N_4762[5]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(spi_data_out_r_39__N_4762[4]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(spi_data_out_r_39__N_4762[3]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(spi_data_out_r_39__N_4762[2]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(spi_data_out_r_39__N_4762[1]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4511[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    LUT4 i12933_2_lut_3_lut (.A(n18666), .B(n18664), .C(n153[0]), .Z(n199[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i12933_2_lut_3_lut.init = 16'h7070;
    LUT4 i13153_2_lut_3_lut (.A(n18666), .B(n18664), .C(n153[1]), .Z(n199[1])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13153_2_lut_3_lut.init = 16'h7070;
    FD1P3AX Cnt_NSL_1780__i11 (.D(n53[11]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780__i11.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1780__i10 (.D(n53[10]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780__i10.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1780__i9 (.D(n53[9]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780__i9.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1780__i8 (.D(n53[8]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780__i8.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1780__i7 (.D(n53[7]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780__i7.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1780__i6 (.D(n53[6]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780__i6.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1780__i5 (.D(n53[5]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780__i5.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1780__i4 (.D(n53[4]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780__i4.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1780__i3 (.D(n53[3]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780__i3.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1780__i2 (.D(n53[2]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780__i2.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1780__i1 (.D(n53[1]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780__i1.GSR = "DISABLED";
    LUT4 i13152_2_lut_3_lut (.A(n18666), .B(n18664), .C(n153[2]), .Z(n199[2])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13152_2_lut_3_lut.init = 16'h7070;
    LUT4 i13151_2_lut_3_lut (.A(n18666), .B(n18664), .C(n153[3]), .Z(n199[3])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13151_2_lut_3_lut.init = 16'h7070;
    FD1S3IX i168_494 (.D(spi_data_out_r_39__N_4848), .CK(clk), .CD(n30185), 
            .Q(spi_data_out_r_39__N_4551)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam i168_494.GSR = "DISABLED";
    FD1P3IX SLO__i43 (.D(SLO[41]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i43.GSR = "DISABLED";
    LUT4 i13150_2_lut_3_lut (.A(n18666), .B(n18664), .C(n153[4]), .Z(n199[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13150_2_lut_3_lut.init = 16'h7070;
    FD1P3IX SLO__i44 (.D(SLO[42]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i44.GSR = "DISABLED";
    FD1P3IX SLO__i45 (.D(SLO[43]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i45.GSR = "DISABLED";
    LUT4 i13149_2_lut_3_lut (.A(n18666), .B(n18664), .C(n153[5]), .Z(n199[5])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13149_2_lut_3_lut.init = 16'h7070;
    FD1P3IX digital_output_r_492 (.D(n28556), .SP(clk_enable_259), .CD(n30185), 
            .CK(clk), .Q(digital_output_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam digital_output_r_492.GSR = "DISABLED";
    LUT4 i13148_2_lut_3_lut (.A(n18666), .B(n18664), .C(n153[6]), .Z(n199[6])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13148_2_lut_3_lut.init = 16'h7070;
    LUT4 i13147_2_lut_3_lut (.A(n18666), .B(n18664), .C(n153[7]), .Z(n199[7])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13147_2_lut_3_lut.init = 16'h7070;
    FD1P3IX SLO__i46 (.D(SLO[44]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i46.GSR = "DISABLED";
    LUT4 mux_158_i1_3_lut (.A(SLO_buf[14]), .B(SLO_buf[4]), .C(n47), .Z(spi_data_out_r_39__N_4762[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i1_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(\quad_homing[0] ), .B(pin_io_c_24), .Z(n25881)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(74[8:17])
    defparam i1_2_lut.init = 16'h8888;
    FD1P3IX mode__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_686), .CD(n30185), 
            .CK(clk), .Q(mode[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i1.GSR = "DISABLED";
    FD1P3IX mode__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_686), .CD(n30185), 
            .CK(clk), .Q(\mode[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i1 (.D(n199[1]), .SP(clk_1MHz_enable_64), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i1.GSR = "DISABLED";
    FD1P3IX Cnt__i2 (.D(n199[2]), .SP(clk_1MHz_enable_64), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i3 (.D(n199[3]), .SP(clk_1MHz_enable_64), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i3.GSR = "DISABLED";
    FD1P3IX Cnt__i4 (.D(n199[4]), .SP(clk_1MHz_enable_64), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i4.GSR = "DISABLED";
    FD1P3IX Cnt__i5 (.D(n199[5]), .SP(clk_1MHz_enable_64), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i5.GSR = "DISABLED";
    FD1P3IX Cnt__i6 (.D(n199[6]), .SP(clk_1MHz_enable_64), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i6.GSR = "DISABLED";
    FD1P3IX Cnt__i7 (.D(n199[7]), .SP(clk_1MHz_enable_64), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i7.GSR = "DISABLED";
    FD1P3AX SLO_buf__i2 (.D(SLO[1]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i2.GSR = "DISABLED";
    FD1P3AX SLO_buf__i3 (.D(SLO[2]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i3.GSR = "DISABLED";
    FD1P3AX SLO_buf__i4 (.D(SLO[3]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i4.GSR = "DISABLED";
    FD1P3AX SLO_buf__i5 (.D(SLO[4]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i5.GSR = "DISABLED";
    FD1P3AX SLO_buf__i6 (.D(SLO[5]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i6.GSR = "DISABLED";
    FD1P3AX SLO_buf__i7 (.D(SLO[6]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i7.GSR = "DISABLED";
    FD1P3AX SLO_buf__i8 (.D(SLO[7]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i8.GSR = "DISABLED";
    FD1P3AX SLO_buf__i9 (.D(SLO[8]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i9.GSR = "DISABLED";
    FD1P3AX SLO_buf__i10 (.D(SLO[9]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i10.GSR = "DISABLED";
    FD1P3AX SLO_buf__i11 (.D(SLO[10]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i11.GSR = "DISABLED";
    FD1P3AX SLO_buf__i12 (.D(SLO[11]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i12.GSR = "DISABLED";
    FD1P3AX SLO_buf__i13 (.D(SLO[12]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i13.GSR = "DISABLED";
    FD1P3AX SLO_buf__i14 (.D(SLO[13]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i14.GSR = "DISABLED";
    FD1P3AX SLO_buf__i15 (.D(SLO[14]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i15.GSR = "DISABLED";
    FD1P3AX SLO_buf__i16 (.D(SLO[15]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i16.GSR = "DISABLED";
    FD1P3AX SLO_buf__i17 (.D(SLO[16]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i17.GSR = "DISABLED";
    FD1P3AX SLO_buf__i18 (.D(SLO[17]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i18.GSR = "DISABLED";
    FD1P3AX SLO_buf__i19 (.D(SLO[18]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i19.GSR = "DISABLED";
    FD1P3AX SLO_buf__i20 (.D(SLO[19]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i20.GSR = "DISABLED";
    FD1P3AX SLO_buf__i21 (.D(SLO[20]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i21.GSR = "DISABLED";
    FD1P3AX SLO_buf__i22 (.D(SLO[21]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i22.GSR = "DISABLED";
    FD1P3AX SLO_buf__i23 (.D(SLO[22]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i23.GSR = "DISABLED";
    FD1P3AX SLO_buf__i24 (.D(SLO[23]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i24.GSR = "DISABLED";
    FD1P3AX SLO_buf__i25 (.D(SLO[24]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i25.GSR = "DISABLED";
    FD1P3AX SLO_buf__i26 (.D(SLO[25]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i26.GSR = "DISABLED";
    FD1P3AX SLO_buf__i27 (.D(SLO[26]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i27.GSR = "DISABLED";
    FD1P3AX SLO_buf__i28 (.D(SLO[27]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i28.GSR = "DISABLED";
    FD1P3AX SLO_buf__i29 (.D(SLO[28]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i29.GSR = "DISABLED";
    FD1P3AX SLO_buf__i30 (.D(SLO[29]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i30.GSR = "DISABLED";
    FD1P3AX SLO_buf__i31 (.D(SLO[30]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i31.GSR = "DISABLED";
    FD1P3AX SLO_buf__i32 (.D(SLO[31]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i32.GSR = "DISABLED";
    FD1P3AX SLO_buf__i33 (.D(SLO[32]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i33.GSR = "DISABLED";
    FD1P3AX SLO_buf__i34 (.D(SLO[33]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i34.GSR = "DISABLED";
    FD1P3AX SLO_buf__i35 (.D(SLO[34]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i35.GSR = "DISABLED";
    FD1P3AX SLO_buf__i36 (.D(SLO[35]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i36.GSR = "DISABLED";
    FD1P3AX SLO_buf__i37 (.D(SLO[36]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i37.GSR = "DISABLED";
    FD1P3AX SLO_buf__i38 (.D(SLO[37]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i38.GSR = "DISABLED";
    FD1P3AX SLO_buf__i39 (.D(SLO[38]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i39.GSR = "DISABLED";
    FD1P3AX SLO_buf__i40 (.D(SLO[39]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i40.GSR = "DISABLED";
    FD1P3AX SLO_buf__i41 (.D(SLO[40]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i41.GSR = "DISABLED";
    FD1P3AX SLO_buf__i42 (.D(SLO[41]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i42.GSR = "DISABLED";
    FD1P3AX SLO_buf__i43 (.D(SLO[42]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i43.GSR = "DISABLED";
    FD1P3AX SLO_buf__i44 (.D(SLO[43]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i44.GSR = "DISABLED";
    FD1P3AX SLO_buf__i45 (.D(SLO[44]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i45.GSR = "DISABLED";
    FD1P3AX SLO_buf__i46 (.D(SLO[45]), .SP(SLO_buf_51__N_4701), .CK(clk), 
            .Q(SLO_buf[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i46.GSR = "DISABLED";
    LUT4 i23966_4_lut (.A(NSL), .B(n30040), .C(n18664), .D(n30003), 
         .Z(NSL_N_4843)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C+(D))))) */ ;
    defparam i23966_4_lut.init = 16'h3b37;
    LUT4 mux_158_i36_3_lut (.A(SLO_buf[9]), .B(SLO_buf[3]), .C(n47), .Z(spi_data_out_r_39__N_4762[35])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i36_3_lut.init = 16'hcaca;
    LUT4 mux_158_i35_3_lut (.A(SLO_buf[8]), .B(SLO_buf[2]), .C(n47), .Z(spi_data_out_r_39__N_4762[34])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i35_3_lut.init = 16'hcaca;
    LUT4 mux_158_i34_3_lut (.A(SLO_buf[7]), .B(SLO_buf[1]), .C(n47), .Z(spi_data_out_r_39__N_4762[33])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i34_3_lut.init = 16'hcaca;
    LUT4 mux_158_i33_3_lut (.A(SLO_buf[6]), .B(SLO_buf[0]), .C(n47), .Z(spi_data_out_r_39__N_4762[32])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i33_3_lut.init = 16'hcaca;
    LUT4 SLO_buf_51__I_142_2_lut (.A(prev_MA_Temp), .B(MA_Temp), .Z(SLO_buf_51__N_4701)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[5:38])
    defparam SLO_buf_51__I_142_2_lut.init = 16'h2222;
    LUT4 mux_158_i16_3_lut (.A(SLO_buf[29]), .B(SLO_buf[19]), .C(n47), 
         .Z(spi_data_out_r_39__N_4762[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i16_3_lut.init = 16'hcaca;
    LUT4 mux_158_i15_3_lut (.A(SLO_buf[28]), .B(SLO_buf[18]), .C(n47), 
         .Z(spi_data_out_r_39__N_4762[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i15_3_lut.init = 16'hcaca;
    LUT4 mux_158_i14_3_lut (.A(SLO_buf[27]), .B(SLO_buf[17]), .C(n47), 
         .Z(spi_data_out_r_39__N_4762[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i14_3_lut.init = 16'hcaca;
    LUT4 mux_158_i13_3_lut (.A(SLO_buf[26]), .B(SLO_buf[16]), .C(n47), 
         .Z(spi_data_out_r_39__N_4762[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i13_3_lut.init = 16'hcaca;
    LUT4 mux_158_i12_3_lut (.A(SLO_buf[25]), .B(SLO_buf[15]), .C(n47), 
         .Z(spi_data_out_r_39__N_4762[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i12_3_lut.init = 16'hcaca;
    LUT4 mux_158_i11_3_lut (.A(SLO_buf[24]), .B(SLO_buf[14]), .C(n47), 
         .Z(spi_data_out_r_39__N_4762[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i11_3_lut.init = 16'hcaca;
    LUT4 mux_158_i10_3_lut (.A(SLO_buf[23]), .B(SLO_buf[13]), .C(n47), 
         .Z(spi_data_out_r_39__N_4762[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i10_3_lut.init = 16'hcaca;
    LUT4 mux_158_i9_3_lut (.A(SLO_buf[22]), .B(SLO_buf[12]), .C(n47), 
         .Z(spi_data_out_r_39__N_4762[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i9_3_lut.init = 16'hcaca;
    LUT4 mux_158_i8_3_lut (.A(SLO_buf[21]), .B(SLO_buf[11]), .C(n47), 
         .Z(spi_data_out_r_39__N_4762[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i8_3_lut.init = 16'hcaca;
    LUT4 mux_158_i7_3_lut (.A(SLO_buf[20]), .B(SLO_buf[10]), .C(n47), 
         .Z(spi_data_out_r_39__N_4762[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i7_3_lut.init = 16'hcaca;
    LUT4 mux_158_i6_3_lut (.A(SLO_buf[19]), .B(SLO_buf[9]), .C(n47), .Z(spi_data_out_r_39__N_4762[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i6_3_lut.init = 16'hcaca;
    LUT4 mux_158_i5_3_lut (.A(SLO_buf[18]), .B(SLO_buf[8]), .C(n47), .Z(spi_data_out_r_39__N_4762[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i5_3_lut.init = 16'hcaca;
    LUT4 mux_158_i4_3_lut (.A(SLO_buf[17]), .B(SLO_buf[7]), .C(n47), .Z(spi_data_out_r_39__N_4762[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i4_3_lut.init = 16'hcaca;
    LUT4 mux_158_i3_3_lut (.A(SLO_buf[16]), .B(SLO_buf[6]), .C(n47), .Z(spi_data_out_r_39__N_4762[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i3_3_lut.init = 16'hcaca;
    LUT4 mux_158_i2_3_lut (.A(SLO_buf[15]), .B(SLO_buf[5]), .C(n47), .Z(spi_data_out_r_39__N_4762[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i2_3_lut.init = 16'hcaca;
    PFUMX MA_Temp_I_157 (.BLUT(n28587), .ALUT(n28588), .C0(n18664), .Z(MA_Temp_N_4830)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;
    LUT4 i24175_4_lut (.A(n30048), .B(n26383), .C(n5), .D(\mode[2] ), 
         .Z(clk_enable_1135)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C)))) */ ;
    defparam i24175_4_lut.init = 16'h0545;
    LUT4 i1_4_lut (.A(mode[1]), .B(mode[0]), .C(Cnt[1]), .D(n4), .Z(n26383)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut.init = 16'h8880;
    CCU2D add_564_9 (.A0(Cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21944), 
          .S0(n153[7]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_9.INIT0 = 16'h5aaa;
    defparam add_564_9.INIT1 = 16'h0000;
    defparam add_564_9.INJECT1_0 = "NO";
    defparam add_564_9.INJECT1_1 = "NO";
    CCU2D add_564_7 (.A0(Cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21943), 
          .COUT(n21944), .S0(n153[5]), .S1(n153[6]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_7.INIT0 = 16'h5aaa;
    defparam add_564_7.INIT1 = 16'h5aaa;
    defparam add_564_7.INJECT1_0 = "NO";
    defparam add_564_7.INJECT1_1 = "NO";
    CCU2D add_564_5 (.A0(Cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21942), 
          .COUT(n21943), .S0(n153[3]), .S1(n153[4]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_5.INIT0 = 16'h5aaa;
    defparam add_564_5.INIT1 = 16'h5aaa;
    defparam add_564_5.INJECT1_0 = "NO";
    defparam add_564_5.INJECT1_1 = "NO";
    CCU2D add_564_3 (.A0(Cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21941), 
          .COUT(n21942), .S0(n153[1]), .S1(n153[2]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_3.INIT0 = 16'h5aaa;
    defparam add_564_3.INIT1 = 16'h5aaa;
    defparam add_564_3.INJECT1_0 = "NO";
    defparam add_564_3.INJECT1_1 = "NO";
    CCU2D add_564_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n21941), 
          .S1(n153[0]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_1.INIT0 = 16'hF000;
    defparam add_564_1.INIT1 = 16'h5555;
    defparam add_564_1.INJECT1_0 = "NO";
    defparam add_564_1.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1780_add_4_13 (.A0(Cnt_NSL[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21933), .S0(n53[11]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780_add_4_13.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1780_add_4_13.INIT1 = 16'h0000;
    defparam Cnt_NSL_1780_add_4_13.INJECT1_0 = "NO";
    defparam Cnt_NSL_1780_add_4_13.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1780_add_4_11 (.A0(Cnt_NSL[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Cnt_NSL[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21932), .COUT(n21933), .S0(n53[9]), .S1(n53[10]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780_add_4_11.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1780_add_4_11.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1780_add_4_11.INJECT1_0 = "NO";
    defparam Cnt_NSL_1780_add_4_11.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1780_add_4_9 (.A0(Cnt_NSL[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Cnt_NSL[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21931), .COUT(n21932), .S0(n53[7]), .S1(n53[8]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780_add_4_9.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1780_add_4_9.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1780_add_4_9.INJECT1_0 = "NO";
    defparam Cnt_NSL_1780_add_4_9.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1780_add_4_7 (.A0(n93[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21930), .COUT(n21931), .S0(n53[5]), .S1(n53[6]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780_add_4_7.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1780_add_4_7.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1780_add_4_7.INJECT1_0 = "NO";
    defparam Cnt_NSL_1780_add_4_7.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1780_add_4_5 (.A0(n93[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21929), .COUT(n21930), .S0(n53[3]), .S1(n53[4]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780_add_4_5.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1780_add_4_5.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1780_add_4_5.INJECT1_0 = "NO";
    defparam Cnt_NSL_1780_add_4_5.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1780_add_4_3 (.A0(n93[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21928), .COUT(n21929), .S0(n53[1]), .S1(n53[2]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780_add_4_3.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1780_add_4_3.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1780_add_4_3.INJECT1_0 = "NO";
    defparam Cnt_NSL_1780_add_4_3.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1780_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n30099), .B1(n30100), .C1(n93[0]), .D1(GND_net), 
          .COUT(n21928), .S1(n53[0]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1780_add_4_1.INIT0 = 16'hF000;
    defparam Cnt_NSL_1780_add_4_1.INIT1 = 16'h8787;
    defparam Cnt_NSL_1780_add_4_1.INJECT1_0 = "NO";
    defparam Cnt_NSL_1780_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_697 (.A(Cnt[7]), .B(Cnt[6]), .Z(n30097)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(109[8:17])
    defparam i1_2_lut_rep_697.init = 16'heeee;
    LUT4 i1_3_lut_rep_668_4_lut (.A(Cnt[7]), .B(Cnt[6]), .C(Cnt[0]), .D(n30202), 
         .Z(n30068)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(109[8:17])
    defparam i1_3_lut_rep_668_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_rep_699 (.A(Cnt_NSL[9]), .B(Cnt_NSL[8]), .C(Cnt_NSL[7]), 
         .Z(n30099)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_rep_699.init = 16'hfefe;
    LUT4 i1_2_lut_rep_640_4_lut (.A(Cnt_NSL[9]), .B(Cnt_NSL[8]), .C(Cnt_NSL[7]), 
         .D(n30100), .Z(n30040)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_rep_640_4_lut.init = 16'hfe00;
    LUT4 i1_2_lut_rep_700 (.A(Cnt_NSL[11]), .B(Cnt_NSL[10]), .Z(n30100)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i1_2_lut_rep_700.init = 16'h8888;
    LUT4 digital_output_r_I_0_547_3_lut (.A(digital_output_r), .B(UC_TXD0_c), 
         .C(OW_ID_N_4805), .Z(OW_ID_N_4804)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[16] 91[59])
    defparam digital_output_r_I_0_547_3_lut.init = 16'hcaca;
    LUT4 i5_4_lut (.A(n9), .B(\uart_slot_en[0] ), .C(n28330), .D(mode[0]), 
         .Z(OW_ID_N_4805)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i5_4_lut.init = 16'h0800;
    LUT4 i23628_2_lut (.A(mode[1]), .B(\uart_slot_en[1] ), .Z(n28330)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23628_2_lut.init = 16'heeee;
    LUT4 i24020_2_lut_rep_615_3_lut_4_lut (.A(Cnt_NSL[11]), .B(Cnt_NSL[10]), 
         .C(resetn_c), .D(n30099), .Z(clk_1MHz_enable_64)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i24020_2_lut_rep_615_3_lut_4_lut.init = 16'h8f0f;
    LUT4 i1_2_lut_rep_802 (.A(Cnt[2]), .B(Cnt[3]), .Z(n30202)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(107[15:23])
    defparam i1_2_lut_rep_802.init = 16'heeee;
    LUT4 i1_3_lut_rep_637_4_lut (.A(Cnt[2]), .B(Cnt[3]), .C(Cnt[1]), .D(Cnt[0]), 
         .Z(n30037)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(107[15:23])
    defparam i1_3_lut_rep_637_4_lut.init = 16'hfeee;
    LUT4 i2978_2_lut_4_lut (.A(mode[1]), .B(mode[0]), .C(\mode[2] ), .D(pin_io_out_29), 
         .Z(\quad_b[2] )) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i2978_2_lut_4_lut.init = 16'h0400;
    LUT4 i2977_2_lut_4_lut (.A(mode[1]), .B(mode[0]), .C(\mode[2] ), .D(pin_io_c_28), 
         .Z(\quad_a[2] )) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i2977_2_lut_4_lut.init = 16'h0400;
    LUT4 i2975_2_lut_3_lut_4_lut (.A(mode[0]), .B(\mode[2] ), .C(pin_io_c_23), 
         .D(mode[1]), .Z(\pin_intrpt[7] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2975_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_2_lut_rep_695_3_lut (.A(mode[0]), .B(\mode[2] ), .C(mode[1]), 
         .Z(n30095)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_rep_695_3_lut.init = 16'hfefe;
    LUT4 i24071_3_lut_4_lut (.A(mode[0]), .B(\mode[2] ), .C(mode[1]), 
         .D(OW_ID_N_4805), .Z(OW_ID_N_4810)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C+(D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i24071_3_lut_4_lut.init = 16'h00ef;
    LUT4 i2974_2_lut_3_lut_4_lut (.A(mode[0]), .B(\mode[2] ), .C(pin_io_c_22), 
         .D(mode[1]), .Z(\pin_intrpt[6] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2974_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2976_2_lut_3_lut_4_lut (.A(mode[0]), .B(\mode[2] ), .C(pin_io_c_24), 
         .D(mode[1]), .Z(\pin_intrpt[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2976_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2959_1_lut_2_lut_3_lut (.A(mode[0]), .B(\mode[2] ), .C(mode[1]), 
         .Z(n7273)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2959_1_lut_2_lut_3_lut.init = 16'h0101;
    LUT4 i2441_2_lut_rep_815 (.A(mode[0]), .B(mode[1]), .Z(n30215)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2441_2_lut_rep_815.init = 16'h8888;
    LUT4 i24074_2_lut_3_lut (.A(mode[0]), .B(mode[1]), .C(\mode[2] ), 
         .Z(ENC_O_N_4812)) /* synthesis lut_function=(!(A (B+(C))+!A (C))) */ ;
    defparam i24074_2_lut_3_lut.init = 16'h0707;
    LUT4 i23931_2_lut_3_lut_4_lut (.A(n30040), .B(resetn_c), .C(n18664), 
         .D(n18666), .Z(clk_1MHz_enable_1)) /* synthesis lut_function=(!(A (C (D))+!A (B+(C (D))))) */ ;
    defparam i23931_2_lut_3_lut_4_lut.init = 16'h0bbb;
    LUT4 i1_2_lut_3_lut (.A(Cnt[5]), .B(n30068), .C(Cnt[4]), .Z(n4)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(133[16:19])
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i23894_1_lut_2_lut_3_lut_4_lut (.A(Cnt[5]), .B(n30068), .C(MA_Temp), 
         .D(n30152), .Z(n28587)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(133[16:19])
    defparam i23894_1_lut_2_lut_3_lut_4_lut.init = 16'he1f0;
    LUT4 i23970_2_lut_rep_710 (.A(MA_Temp), .B(clk_1MHz), .Z(n30110)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i23970_2_lut_rep_710.init = 16'h7777;
    LUT4 i23940_2_lut_3_lut_4_lut (.A(MA_Temp), .B(clk_1MHz), .C(n5), 
         .D(prev_MA), .Z(n12391)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i23940_2_lut_3_lut_4_lut.init = 16'h0007;
    LUT4 i1_2_lut_rep_648_3_lut (.A(MA_Temp), .B(clk_1MHz), .C(prev_MA), 
         .Z(n30048)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i1_2_lut_rep_648_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut (.A(mode[1]), .B(\mode[2] ), .C(mode[0]), .Z(n5)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_3_lut.init = 16'hfbfb;
    FD1P3AX NSL_484 (.D(NSL_N_4843), .SP(clk_1MHz_enable_66), .CK(clk_1MHz), 
            .Q(NSL)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam NSL_484.GSR = "DISABLED";
    FD1P3IX SLO__i24 (.D(SLO[22]), .SP(clk_enable_1135), .CD(n12391), 
            .CK(clk), .Q(SLO[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i24.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_849 (.A(n30097), .B(n24971), .C(n30215), .D(\mode[2] ), 
         .Z(n18666)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i1_4_lut_adj_849.init = 16'hffef;
    LUT4 i1_3_lut_adj_850 (.A(Cnt[5]), .B(n30037), .C(Cnt[4]), .Z(n24971)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_850.init = 16'h8080;
    LUT4 i1_4_lut_adj_851 (.A(n30097), .B(n18578), .C(Cnt[5]), .D(n5), 
         .Z(n18664)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_851.init = 16'hfffe;
    LUT4 i13288_2_lut_rep_752 (.A(Cnt[4]), .B(Cnt[1]), .Z(n30152)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13288_2_lut_rep_752.init = 16'h8888;
    LUT4 i23616_2_lut_3_lut (.A(Cnt[4]), .B(Cnt[1]), .C(Cnt[5]), .Z(n28318)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i23616_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_603_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(n30068), 
         .D(Cnt[5]), .Z(n30003)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_rep_603_3_lut_4_lut.init = 16'hfff7;
    
endmodule
//
// Verilog Description of module \quad_decoder(DEV_ID=5) 
//

module \quad_decoder(DEV_ID=5)  (quad_homing, clk, clk_enable_388, n30185, 
            \spi_data_r[0] , quad_count, \quad_b[5] , \spi_data_out_r_39__N_2109[0] , 
            \spi_data_out_r_39__N_2258[0] , quad_buffer, \pin_intrpt[17] , 
            GND_net, clk_enable_315, \quad_a[5] , spi_data_out_r_39__N_2149, 
            spi_data_out_r_39__N_2338, quad_set_valid_N_2333, \spi_data_r[31] , 
            \spi_data_r[30] , \spi_data_r[29] , \spi_data_r[28] , \spi_data_r[27] , 
            \spi_data_r[26] , \spi_data_r[25] , \spi_data_r[24] , \spi_data_r[23] , 
            \spi_data_r[22] , \spi_data_r[21] , \spi_data_r[20] , \spi_data_r[19] , 
            \spi_data_r[18] , \spi_data_r[17] , \spi_data_r[16] , \spi_data_r[15] , 
            \spi_data_r[14] , \spi_data_r[13] , \spi_data_r[12] , \spi_data_r[11] , 
            \spi_data_r[10] , \spi_data_r[9] , \spi_data_r[8] , \spi_data_r[7] , 
            \spi_data_r[6] , \spi_data_r[5] , \spi_data_r[4] , \spi_data_r[3] , 
            \spi_data_r[2] , \spi_data_r[1] , \spi_data_out_r_39__N_2109[31] , 
            \spi_data_out_r_39__N_2258[31] , \spi_data_out_r_39__N_2109[30] , 
            \spi_data_out_r_39__N_2258[30] , \spi_data_out_r_39__N_2109[29] , 
            \spi_data_out_r_39__N_2258[29] , \spi_data_out_r_39__N_2109[28] , 
            \spi_data_out_r_39__N_2258[28] , \spi_data_out_r_39__N_2109[27] , 
            \spi_data_out_r_39__N_2258[27] , \spi_data_out_r_39__N_2109[26] , 
            \spi_data_out_r_39__N_2258[26] , \spi_data_out_r_39__N_2109[25] , 
            \spi_data_out_r_39__N_2258[25] , \spi_data_out_r_39__N_2109[24] , 
            \spi_data_out_r_39__N_2258[24] , \spi_data_out_r_39__N_2109[23] , 
            \spi_data_out_r_39__N_2258[23] , \spi_data_out_r_39__N_2109[22] , 
            \spi_data_out_r_39__N_2258[22] , \spi_data_out_r_39__N_2109[21] , 
            \spi_data_out_r_39__N_2258[21] , \spi_data_out_r_39__N_2109[20] , 
            \spi_data_out_r_39__N_2258[20] , \spi_data_out_r_39__N_2109[19] , 
            \spi_data_out_r_39__N_2258[19] , \spi_data_out_r_39__N_2109[18] , 
            \spi_data_out_r_39__N_2258[18] , \spi_data_out_r_39__N_2109[17] , 
            \spi_data_out_r_39__N_2258[17] , \spi_data_out_r_39__N_2109[16] , 
            \spi_data_out_r_39__N_2258[16] , \spi_data_out_r_39__N_2109[15] , 
            \spi_data_out_r_39__N_2258[15] , \spi_data_out_r_39__N_2109[14] , 
            \spi_data_out_r_39__N_2258[14] , \spi_data_out_r_39__N_2109[13] , 
            \spi_data_out_r_39__N_2258[13] , \spi_data_out_r_39__N_2109[12] , 
            \spi_data_out_r_39__N_2258[12] , \spi_data_out_r_39__N_2109[11] , 
            \spi_data_out_r_39__N_2258[11] , \spi_data_out_r_39__N_2109[10] , 
            \spi_data_out_r_39__N_2258[10] , \spi_data_out_r_39__N_2109[9] , 
            \spi_data_out_r_39__N_2258[9] , \spi_data_out_r_39__N_2109[8] , 
            \spi_data_out_r_39__N_2258[8] , \spi_data_out_r_39__N_2109[7] , 
            \spi_data_out_r_39__N_2258[7] , \spi_data_out_r_39__N_2109[6] , 
            \spi_data_out_r_39__N_2258[6] , \spi_data_out_r_39__N_2109[5] , 
            \spi_data_out_r_39__N_2258[5] , \spi_data_out_r_39__N_2109[4] , 
            \spi_data_out_r_39__N_2258[4] , \spi_data_out_r_39__N_2109[3] , 
            \spi_data_out_r_39__N_2258[3] , \spi_data_out_r_39__N_2109[2] , 
            \spi_data_out_r_39__N_2258[2] , \spi_data_out_r_39__N_2109[1] , 
            \spi_data_out_r_39__N_2258[1] , resetn_c, n1) /* synthesis syn_module_defined=1 */ ;
    output [1:0]quad_homing;
    input clk;
    input clk_enable_388;
    input n30185;
    input \spi_data_r[0] ;
    output [31:0]quad_count;
    input \quad_b[5] ;
    output \spi_data_out_r_39__N_2109[0] ;
    input \spi_data_out_r_39__N_2258[0] ;
    output [31:0]quad_buffer;
    input \pin_intrpt[17] ;
    input GND_net;
    input clk_enable_315;
    input \quad_a[5] ;
    output spi_data_out_r_39__N_2149;
    input spi_data_out_r_39__N_2338;
    input quad_set_valid_N_2333;
    input \spi_data_r[31] ;
    input \spi_data_r[30] ;
    input \spi_data_r[29] ;
    input \spi_data_r[28] ;
    input \spi_data_r[27] ;
    input \spi_data_r[26] ;
    input \spi_data_r[25] ;
    input \spi_data_r[24] ;
    input \spi_data_r[23] ;
    input \spi_data_r[22] ;
    input \spi_data_r[21] ;
    input \spi_data_r[20] ;
    input \spi_data_r[19] ;
    input \spi_data_r[18] ;
    input \spi_data_r[17] ;
    input \spi_data_r[16] ;
    input \spi_data_r[15] ;
    input \spi_data_r[14] ;
    input \spi_data_r[13] ;
    input \spi_data_r[12] ;
    input \spi_data_r[11] ;
    input \spi_data_r[10] ;
    input \spi_data_r[9] ;
    input \spi_data_r[8] ;
    input \spi_data_r[7] ;
    input \spi_data_r[6] ;
    input \spi_data_r[5] ;
    input \spi_data_r[4] ;
    input \spi_data_r[3] ;
    input \spi_data_r[2] ;
    input \spi_data_r[1] ;
    output \spi_data_out_r_39__N_2109[31] ;
    input \spi_data_out_r_39__N_2258[31] ;
    output \spi_data_out_r_39__N_2109[30] ;
    input \spi_data_out_r_39__N_2258[30] ;
    output \spi_data_out_r_39__N_2109[29] ;
    input \spi_data_out_r_39__N_2258[29] ;
    output \spi_data_out_r_39__N_2109[28] ;
    input \spi_data_out_r_39__N_2258[28] ;
    output \spi_data_out_r_39__N_2109[27] ;
    input \spi_data_out_r_39__N_2258[27] ;
    output \spi_data_out_r_39__N_2109[26] ;
    input \spi_data_out_r_39__N_2258[26] ;
    output \spi_data_out_r_39__N_2109[25] ;
    input \spi_data_out_r_39__N_2258[25] ;
    output \spi_data_out_r_39__N_2109[24] ;
    input \spi_data_out_r_39__N_2258[24] ;
    output \spi_data_out_r_39__N_2109[23] ;
    input \spi_data_out_r_39__N_2258[23] ;
    output \spi_data_out_r_39__N_2109[22] ;
    input \spi_data_out_r_39__N_2258[22] ;
    output \spi_data_out_r_39__N_2109[21] ;
    input \spi_data_out_r_39__N_2258[21] ;
    output \spi_data_out_r_39__N_2109[20] ;
    input \spi_data_out_r_39__N_2258[20] ;
    output \spi_data_out_r_39__N_2109[19] ;
    input \spi_data_out_r_39__N_2258[19] ;
    output \spi_data_out_r_39__N_2109[18] ;
    input \spi_data_out_r_39__N_2258[18] ;
    output \spi_data_out_r_39__N_2109[17] ;
    input \spi_data_out_r_39__N_2258[17] ;
    output \spi_data_out_r_39__N_2109[16] ;
    input \spi_data_out_r_39__N_2258[16] ;
    output \spi_data_out_r_39__N_2109[15] ;
    input \spi_data_out_r_39__N_2258[15] ;
    output \spi_data_out_r_39__N_2109[14] ;
    input \spi_data_out_r_39__N_2258[14] ;
    output \spi_data_out_r_39__N_2109[13] ;
    input \spi_data_out_r_39__N_2258[13] ;
    output \spi_data_out_r_39__N_2109[12] ;
    input \spi_data_out_r_39__N_2258[12] ;
    output \spi_data_out_r_39__N_2109[11] ;
    input \spi_data_out_r_39__N_2258[11] ;
    output \spi_data_out_r_39__N_2109[10] ;
    input \spi_data_out_r_39__N_2258[10] ;
    output \spi_data_out_r_39__N_2109[9] ;
    input \spi_data_out_r_39__N_2258[9] ;
    output \spi_data_out_r_39__N_2109[8] ;
    input \spi_data_out_r_39__N_2258[8] ;
    output \spi_data_out_r_39__N_2109[7] ;
    input \spi_data_out_r_39__N_2258[7] ;
    output \spi_data_out_r_39__N_2109[6] ;
    input \spi_data_out_r_39__N_2258[6] ;
    output \spi_data_out_r_39__N_2109[5] ;
    input \spi_data_out_r_39__N_2258[5] ;
    output \spi_data_out_r_39__N_2109[4] ;
    input \spi_data_out_r_39__N_2258[4] ;
    output \spi_data_out_r_39__N_2109[3] ;
    input \spi_data_out_r_39__N_2258[3] ;
    output \spi_data_out_r_39__N_2109[2] ;
    input \spi_data_out_r_39__N_2258[2] ;
    output \spi_data_out_r_39__N_2109[1] ;
    input \spi_data_out_r_39__N_2258[1] ;
    input resetn_c;
    input n1;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire \pin_intrpt[17]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[17] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    
    wire clk_enable_385, n7953;
    wire [2:0]quad_b_delayed;   // c:/s_links/sources/quad_decoder.v(35[19:33])
    wire [2:0]quad_a_delayed;   // c:/s_links/sources/quad_decoder.v(34[20:34])
    
    wire n21844;
    wire [31:0]quad_set;   // c:/s_links/sources/quad_decoder.v(39[31:39])
    
    wire quad_set_valid, n8807, n8809, n8811, n8813, n8815, n8817, 
        n8819, n8821, n8823, n8825, n8827, n8829, n8831, n8833, 
        n8835, n8837, n8839, n8841, n8843, n8845, n8847, n8849, 
        n8851, n8853, n8855, n8857, n8859, n8861, n8863, n8865, 
        n8867, n6, count_dir, n21859;
    wire [31:0]n3930;
    
    wire n21858, n21857, n21856, n21855, n21854, n21853, n21852, 
        n5717, n21851, n21850, n21849, n21848, n21847, n21846, 
        n21845;
    
    FD1P3IX quad_homing__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_388), .CD(n30185), 
            .CK(clk), .Q(quad_homing[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(62[8] 69[4])
    defparam quad_homing__i0.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i0 (.D(n7953), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i0.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i0 (.D(\quad_b[5] ), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_2258[0] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX quad_buffer_i0 (.D(quad_count[0]), .CK(\pin_intrpt[17] ), .Q(quad_buffer[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i0.GSR = "DISABLED";
    CCU2D add_1385_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quad_a_delayed[2]), .B1(quad_b_delayed[1]), .C1(quad_b_delayed[2]), 
          .D1(quad_a_delayed[1]), .COUT(n21844));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_1.INIT0 = 16'hF000;
    defparam add_1385_1.INIT1 = 16'h0990;
    defparam add_1385_1.INJECT1_0 = "NO";
    defparam add_1385_1.INJECT1_1 = "NO";
    FD1P3IX quad_set__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i0.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i0 (.D(\quad_a[5] ), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i0.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i2 (.D(quad_a_delayed[1]), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i2.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i1 (.D(quad_a_delayed[0]), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i1.GSR = "DISABLED";
    FD1S3IX i39_391 (.D(spi_data_out_r_39__N_2338), .CK(clk), .CD(n30185), 
            .Q(spi_data_out_r_39__N_2149)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam i39_391.GSR = "DISABLED";
    FD1S3IX quad_set_valid_388 (.D(quad_set_valid_N_2333), .CK(clk), .CD(n30185), 
            .Q(quad_set_valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set_valid_388.GSR = "DISABLED";
    FD1P3IX quad_set__i31 (.D(\spi_data_r[31] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i31.GSR = "DISABLED";
    FD1P3IX quad_set__i30 (.D(\spi_data_r[30] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i30.GSR = "DISABLED";
    FD1P3IX quad_set__i29 (.D(\spi_data_r[29] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i29.GSR = "DISABLED";
    FD1P3IX quad_set__i28 (.D(\spi_data_r[28] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i28.GSR = "DISABLED";
    FD1P3IX quad_set__i27 (.D(\spi_data_r[27] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i27.GSR = "DISABLED";
    FD1P3IX quad_set__i26 (.D(\spi_data_r[26] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i26.GSR = "DISABLED";
    FD1P3IX quad_set__i25 (.D(\spi_data_r[25] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i25.GSR = "DISABLED";
    FD1P3IX quad_set__i24 (.D(\spi_data_r[24] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i24.GSR = "DISABLED";
    FD1P3IX quad_set__i23 (.D(\spi_data_r[23] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i23.GSR = "DISABLED";
    FD1P3IX quad_set__i22 (.D(\spi_data_r[22] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i22.GSR = "DISABLED";
    FD1P3IX quad_set__i21 (.D(\spi_data_r[21] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i21.GSR = "DISABLED";
    FD1P3IX quad_set__i20 (.D(\spi_data_r[20] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i20.GSR = "DISABLED";
    FD1P3IX quad_set__i19 (.D(\spi_data_r[19] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i19.GSR = "DISABLED";
    FD1P3IX quad_set__i18 (.D(\spi_data_r[18] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i18.GSR = "DISABLED";
    FD1P3IX quad_set__i17 (.D(\spi_data_r[17] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i17.GSR = "DISABLED";
    FD1P3IX quad_set__i16 (.D(\spi_data_r[16] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i16.GSR = "DISABLED";
    FD1P3IX quad_set__i15 (.D(\spi_data_r[15] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i15.GSR = "DISABLED";
    FD1P3IX quad_set__i14 (.D(\spi_data_r[14] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i14.GSR = "DISABLED";
    FD1P3IX quad_set__i13 (.D(\spi_data_r[13] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i13.GSR = "DISABLED";
    FD1P3IX quad_set__i12 (.D(\spi_data_r[12] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i12.GSR = "DISABLED";
    FD1P3IX quad_set__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i11.GSR = "DISABLED";
    FD1P3IX quad_set__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i10.GSR = "DISABLED";
    FD1P3IX quad_set__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i9.GSR = "DISABLED";
    FD1P3IX quad_set__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i8.GSR = "DISABLED";
    FD1P3IX quad_set__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i7.GSR = "DISABLED";
    FD1P3IX quad_set__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i6.GSR = "DISABLED";
    FD1P3IX quad_set__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i5.GSR = "DISABLED";
    FD1P3IX quad_set__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i4.GSR = "DISABLED";
    FD1P3IX quad_set__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i3.GSR = "DISABLED";
    FD1P3IX quad_set__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i2.GSR = "DISABLED";
    FD1P3IX quad_set__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_315), .CD(n30185), 
            .CK(clk), .Q(quad_set[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i1.GSR = "DISABLED";
    FD1S3AX quad_buffer_i31 (.D(quad_count[31]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i31.GSR = "DISABLED";
    FD1S3AX quad_buffer_i30 (.D(quad_count[30]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i30.GSR = "DISABLED";
    FD1S3AX quad_buffer_i29 (.D(quad_count[29]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i29.GSR = "DISABLED";
    FD1S3AX quad_buffer_i28 (.D(quad_count[28]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i28.GSR = "DISABLED";
    FD1S3AX quad_buffer_i27 (.D(quad_count[27]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i27.GSR = "DISABLED";
    FD1S3AX quad_buffer_i26 (.D(quad_count[26]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i26.GSR = "DISABLED";
    FD1S3AX quad_buffer_i25 (.D(quad_count[25]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i25.GSR = "DISABLED";
    FD1S3AX quad_buffer_i24 (.D(quad_count[24]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i24.GSR = "DISABLED";
    FD1S3AX quad_buffer_i23 (.D(quad_count[23]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i23.GSR = "DISABLED";
    FD1S3AX quad_buffer_i22 (.D(quad_count[22]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i22.GSR = "DISABLED";
    FD1S3AX quad_buffer_i21 (.D(quad_count[21]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i21.GSR = "DISABLED";
    FD1S3AX quad_buffer_i20 (.D(quad_count[20]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i20.GSR = "DISABLED";
    FD1S3AX quad_buffer_i19 (.D(quad_count[19]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i19.GSR = "DISABLED";
    FD1S3AX quad_buffer_i18 (.D(quad_count[18]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i18.GSR = "DISABLED";
    FD1S3AX quad_buffer_i17 (.D(quad_count[17]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i17.GSR = "DISABLED";
    FD1S3AX quad_buffer_i16 (.D(quad_count[16]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i16.GSR = "DISABLED";
    FD1S3AX quad_buffer_i15 (.D(quad_count[15]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i15.GSR = "DISABLED";
    FD1S3AX quad_buffer_i14 (.D(quad_count[14]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i14.GSR = "DISABLED";
    FD1S3AX quad_buffer_i13 (.D(quad_count[13]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i13.GSR = "DISABLED";
    FD1S3AX quad_buffer_i12 (.D(quad_count[12]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i12.GSR = "DISABLED";
    FD1S3AX quad_buffer_i11 (.D(quad_count[11]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i11.GSR = "DISABLED";
    FD1S3AX quad_buffer_i10 (.D(quad_count[10]), .CK(\pin_intrpt[17] ), 
            .Q(quad_buffer[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i10.GSR = "DISABLED";
    FD1S3AX quad_buffer_i9 (.D(quad_count[9]), .CK(\pin_intrpt[17] ), .Q(quad_buffer[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i9.GSR = "DISABLED";
    FD1S3AX quad_buffer_i8 (.D(quad_count[8]), .CK(\pin_intrpt[17] ), .Q(quad_buffer[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i8.GSR = "DISABLED";
    FD1S3AX quad_buffer_i7 (.D(quad_count[7]), .CK(\pin_intrpt[17] ), .Q(quad_buffer[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i7.GSR = "DISABLED";
    FD1S3AX quad_buffer_i6 (.D(quad_count[6]), .CK(\pin_intrpt[17] ), .Q(quad_buffer[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i6.GSR = "DISABLED";
    FD1S3AX quad_buffer_i5 (.D(quad_count[5]), .CK(\pin_intrpt[17] ), .Q(quad_buffer[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i5.GSR = "DISABLED";
    FD1S3AX quad_buffer_i4 (.D(quad_count[4]), .CK(\pin_intrpt[17] ), .Q(quad_buffer[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i4.GSR = "DISABLED";
    FD1S3AX quad_buffer_i3 (.D(quad_count[3]), .CK(\pin_intrpt[17] ), .Q(quad_buffer[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i3.GSR = "DISABLED";
    FD1S3AX quad_buffer_i2 (.D(quad_count[2]), .CK(\pin_intrpt[17] ), .Q(quad_buffer[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i2.GSR = "DISABLED";
    FD1S3AX quad_buffer_i1 (.D(quad_count[1]), .CK(\pin_intrpt[17] ), .Q(quad_buffer[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_2258[31] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i31 (.D(\spi_data_out_r_39__N_2258[30] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i30 (.D(\spi_data_out_r_39__N_2258[29] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i29 (.D(\spi_data_out_r_39__N_2258[28] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i28 (.D(\spi_data_out_r_39__N_2258[27] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i27 (.D(\spi_data_out_r_39__N_2258[26] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i26 (.D(\spi_data_out_r_39__N_2258[25] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i25 (.D(\spi_data_out_r_39__N_2258[24] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i24 (.D(\spi_data_out_r_39__N_2258[23] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i23 (.D(\spi_data_out_r_39__N_2258[22] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i22 (.D(\spi_data_out_r_39__N_2258[21] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i21 (.D(\spi_data_out_r_39__N_2258[20] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i20 (.D(\spi_data_out_r_39__N_2258[19] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i19 (.D(\spi_data_out_r_39__N_2258[18] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i18 (.D(\spi_data_out_r_39__N_2258[17] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i17 (.D(\spi_data_out_r_39__N_2258[16] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i16 (.D(\spi_data_out_r_39__N_2258[15] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_2258[14] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_2258[13] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_2258[12] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_2258[11] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_2258[10] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_2258[9] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_2258[8] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_2258[7] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_2258[6] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_2258[5] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_2258[4] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_2258[3] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_2258[2] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_2258[1] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2109[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i2 (.D(quad_b_delayed[1]), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i2.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i1 (.D(quad_b_delayed[0]), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i1.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i31 (.D(n8807), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i31.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i30 (.D(n8809), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i30.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i29 (.D(n8811), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i29.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i28 (.D(n8813), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i28.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i27 (.D(n8815), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i27.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i26 (.D(n8817), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i26.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i25 (.D(n8819), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i25.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i24 (.D(n8821), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i24.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i23 (.D(n8823), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i23.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i22 (.D(n8825), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i22.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i21 (.D(n8827), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i21.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i20 (.D(n8829), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i20.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i19 (.D(n8831), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i19.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i18 (.D(n8833), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i18.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i17 (.D(n8835), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i17.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i16 (.D(n8837), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i16.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i15 (.D(n8839), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i15.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i14 (.D(n8841), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i14.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i13 (.D(n8843), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i13.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i12 (.D(n8845), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i12.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i11 (.D(n8847), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i11.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i10 (.D(n8849), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i10.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i9 (.D(n8851), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i9.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i8 (.D(n8853), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i8.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i7 (.D(n8855), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i7.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i6 (.D(n8857), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i6.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i5 (.D(n8859), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i5.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i4 (.D(n8861), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i4.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i3 (.D(n8863), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i3.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i2 (.D(n8865), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i1 (.D(n8867), .SP(clk_enable_385), .CK(clk), 
            .Q(quad_count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i1.GSR = "DISABLED";
    FD1P3IX quad_homing__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_388), .CD(n30185), 
            .CK(clk), .Q(quad_homing[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(62[8] 69[4])
    defparam quad_homing__i1.GSR = "DISABLED";
    LUT4 i2_2_lut (.A(quad_b_delayed[1]), .B(quad_a_delayed[2]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(96[19:96])
    defparam i2_2_lut.init = 16'h6666;
    LUT4 i1_2_lut (.A(quad_a_delayed[1]), .B(quad_b_delayed[2]), .Z(count_dir)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(96[19:96])
    defparam i1_2_lut.init = 16'h6666;
    CCU2D add_1385_33 (.A0(quad_count[30]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[31]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21859), .S0(n3930[30]), .S1(n3930[31]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_33.INIT0 = 16'h5569;
    defparam add_1385_33.INIT1 = 16'h5569;
    defparam add_1385_33.INJECT1_0 = "NO";
    defparam add_1385_33.INJECT1_1 = "NO";
    CCU2D add_1385_31 (.A0(quad_count[28]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[29]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21858), .COUT(n21859), .S0(n3930[28]), .S1(n3930[29]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_31.INIT0 = 16'h5569;
    defparam add_1385_31.INIT1 = 16'h5569;
    defparam add_1385_31.INJECT1_0 = "NO";
    defparam add_1385_31.INJECT1_1 = "NO";
    CCU2D add_1385_29 (.A0(quad_count[26]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[27]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21857), .COUT(n21858), .S0(n3930[26]), .S1(n3930[27]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_29.INIT0 = 16'h5569;
    defparam add_1385_29.INIT1 = 16'h5569;
    defparam add_1385_29.INJECT1_0 = "NO";
    defparam add_1385_29.INJECT1_1 = "NO";
    LUT4 i24187_2_lut (.A(resetn_c), .B(quad_homing[1]), .Z(clk_enable_385)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i24187_2_lut.init = 16'h7777;
    CCU2D add_1385_27 (.A0(quad_count[24]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[25]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21856), .COUT(n21857), .S0(n3930[24]), .S1(n3930[25]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_27.INIT0 = 16'h5569;
    defparam add_1385_27.INIT1 = 16'h5569;
    defparam add_1385_27.INJECT1_0 = "NO";
    defparam add_1385_27.INJECT1_1 = "NO";
    CCU2D add_1385_25 (.A0(quad_count[22]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[23]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21855), .COUT(n21856), .S0(n3930[22]), .S1(n3930[23]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_25.INIT0 = 16'h5569;
    defparam add_1385_25.INIT1 = 16'h5569;
    defparam add_1385_25.INJECT1_0 = "NO";
    defparam add_1385_25.INJECT1_1 = "NO";
    CCU2D add_1385_23 (.A0(quad_count[20]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[21]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21854), .COUT(n21855), .S0(n3930[20]), .S1(n3930[21]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_23.INIT0 = 16'h5569;
    defparam add_1385_23.INIT1 = 16'h5569;
    defparam add_1385_23.INJECT1_0 = "NO";
    defparam add_1385_23.INJECT1_1 = "NO";
    CCU2D add_1385_21 (.A0(quad_count[18]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[19]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21853), .COUT(n21854), .S0(n3930[18]), .S1(n3930[19]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_21.INIT0 = 16'h5569;
    defparam add_1385_21.INIT1 = 16'h5569;
    defparam add_1385_21.INJECT1_0 = "NO";
    defparam add_1385_21.INJECT1_1 = "NO";
    CCU2D add_1385_19 (.A0(quad_count[16]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[17]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21852), .COUT(n21853), .S0(n3930[16]), .S1(n3930[17]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_19.INIT0 = 16'h5569;
    defparam add_1385_19.INIT1 = 16'h5569;
    defparam add_1385_19.INJECT1_0 = "NO";
    defparam add_1385_19.INJECT1_1 = "NO";
    LUT4 i3631_4_lut (.A(n3930[0]), .B(quad_set[0]), .C(n5717), .D(n1), 
         .Z(n7953)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i3631_4_lut.init = 16'hc0ca;
    CCU2D add_1385_17 (.A0(quad_count[14]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[15]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21851), .COUT(n21852), .S0(n3930[14]), .S1(n3930[15]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_17.INIT0 = 16'h5569;
    defparam add_1385_17.INIT1 = 16'h5569;
    defparam add_1385_17.INJECT1_0 = "NO";
    defparam add_1385_17.INJECT1_1 = "NO";
    CCU2D add_1385_15 (.A0(quad_count[12]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[13]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21850), .COUT(n21851), .S0(n3930[12]), .S1(n3930[13]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_15.INIT0 = 16'h5569;
    defparam add_1385_15.INIT1 = 16'h5569;
    defparam add_1385_15.INJECT1_0 = "NO";
    defparam add_1385_15.INJECT1_1 = "NO";
    CCU2D add_1385_13 (.A0(quad_count[10]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[11]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21849), .COUT(n21850), .S0(n3930[10]), .S1(n3930[11]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_13.INIT0 = 16'h5569;
    defparam add_1385_13.INIT1 = 16'h5569;
    defparam add_1385_13.INJECT1_0 = "NO";
    defparam add_1385_13.INJECT1_1 = "NO";
    CCU2D add_1385_11 (.A0(quad_count[8]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[9]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21848), .COUT(n21849), .S0(n3930[8]), .S1(n3930[9]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_11.INIT0 = 16'h5569;
    defparam add_1385_11.INIT1 = 16'h5569;
    defparam add_1385_11.INJECT1_0 = "NO";
    defparam add_1385_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(quad_homing[0]), .B(quad_homing[1]), .C(quad_set_valid), 
         .D(resetn_c), .Z(n5717)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut.init = 16'h1000;
    CCU2D add_1385_9 (.A0(quad_count[6]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[7]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21847), .COUT(n21848), .S0(n3930[6]), .S1(n3930[7]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_9.INIT0 = 16'h5569;
    defparam add_1385_9.INIT1 = 16'h5569;
    defparam add_1385_9.INJECT1_0 = "NO";
    defparam add_1385_9.INJECT1_1 = "NO";
    CCU2D add_1385_7 (.A0(quad_count[4]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[5]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21846), .COUT(n21847), .S0(n3930[4]), .S1(n3930[5]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_7.INIT0 = 16'h5569;
    defparam add_1385_7.INIT1 = 16'h5569;
    defparam add_1385_7.INJECT1_0 = "NO";
    defparam add_1385_7.INJECT1_1 = "NO";
    CCU2D add_1385_5 (.A0(quad_count[2]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[3]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21845), .COUT(n21846), .S0(n3930[2]), .S1(n3930[3]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_5.INIT0 = 16'h5569;
    defparam add_1385_5.INIT1 = 16'h5569;
    defparam add_1385_5.INJECT1_0 = "NO";
    defparam add_1385_5.INJECT1_1 = "NO";
    CCU2D add_1385_3 (.A0(quad_count[0]), .B0(count_dir), .C0(n6), .D0(count_dir), 
          .A1(quad_count[1]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21844), .COUT(n21845), .S0(n3930[0]), .S1(n3930[1]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1385_3.INIT0 = 16'h5665;
    defparam add_1385_3.INIT1 = 16'h5569;
    defparam add_1385_3.INJECT1_0 = "NO";
    defparam add_1385_3.INJECT1_1 = "NO";
    LUT4 i4483_4_lut (.A(n3930[31]), .B(quad_set[31]), .C(n5717), .D(n1), 
         .Z(n8807)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4483_4_lut.init = 16'hc0ca;
    LUT4 i4485_4_lut (.A(n3930[30]), .B(quad_set[30]), .C(n5717), .D(n1), 
         .Z(n8809)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4485_4_lut.init = 16'hc0ca;
    LUT4 i4487_4_lut (.A(n3930[29]), .B(quad_set[29]), .C(n5717), .D(n1), 
         .Z(n8811)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4487_4_lut.init = 16'hc0ca;
    LUT4 i4489_4_lut (.A(n3930[28]), .B(quad_set[28]), .C(n5717), .D(n1), 
         .Z(n8813)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4489_4_lut.init = 16'hc0ca;
    LUT4 i4491_4_lut (.A(n3930[27]), .B(quad_set[27]), .C(n5717), .D(n1), 
         .Z(n8815)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4491_4_lut.init = 16'hc0ca;
    LUT4 i4493_4_lut (.A(n3930[26]), .B(quad_set[26]), .C(n5717), .D(n1), 
         .Z(n8817)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4493_4_lut.init = 16'hc0ca;
    LUT4 i4495_4_lut (.A(n3930[25]), .B(quad_set[25]), .C(n5717), .D(n1), 
         .Z(n8819)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4495_4_lut.init = 16'hc0ca;
    LUT4 i4497_4_lut (.A(n3930[24]), .B(quad_set[24]), .C(n5717), .D(n1), 
         .Z(n8821)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4497_4_lut.init = 16'hc0ca;
    LUT4 i4499_4_lut (.A(n3930[23]), .B(quad_set[23]), .C(n5717), .D(n1), 
         .Z(n8823)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4499_4_lut.init = 16'hc0ca;
    LUT4 i4501_4_lut (.A(n3930[22]), .B(quad_set[22]), .C(n5717), .D(n1), 
         .Z(n8825)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4501_4_lut.init = 16'hc0ca;
    LUT4 i4503_4_lut (.A(n3930[21]), .B(quad_set[21]), .C(n5717), .D(n1), 
         .Z(n8827)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4503_4_lut.init = 16'hc0ca;
    LUT4 i4505_4_lut (.A(n3930[20]), .B(quad_set[20]), .C(n5717), .D(n1), 
         .Z(n8829)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4505_4_lut.init = 16'hc0ca;
    LUT4 i4507_4_lut (.A(n3930[19]), .B(quad_set[19]), .C(n5717), .D(n1), 
         .Z(n8831)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4507_4_lut.init = 16'hc0ca;
    LUT4 i4509_4_lut (.A(n3930[18]), .B(quad_set[18]), .C(n5717), .D(n1), 
         .Z(n8833)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4509_4_lut.init = 16'hc0ca;
    LUT4 i4511_4_lut (.A(n3930[17]), .B(quad_set[17]), .C(n5717), .D(n1), 
         .Z(n8835)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4511_4_lut.init = 16'hc0ca;
    LUT4 i4513_4_lut (.A(n3930[16]), .B(quad_set[16]), .C(n5717), .D(n1), 
         .Z(n8837)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4513_4_lut.init = 16'hc0ca;
    LUT4 i4515_4_lut (.A(n3930[15]), .B(quad_set[15]), .C(n5717), .D(n1), 
         .Z(n8839)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4515_4_lut.init = 16'hc0ca;
    LUT4 i4517_4_lut (.A(n3930[14]), .B(quad_set[14]), .C(n5717), .D(n1), 
         .Z(n8841)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4517_4_lut.init = 16'hc0ca;
    LUT4 i4519_4_lut (.A(n3930[13]), .B(quad_set[13]), .C(n5717), .D(n1), 
         .Z(n8843)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4519_4_lut.init = 16'hc0ca;
    LUT4 i4521_4_lut (.A(n3930[12]), .B(quad_set[12]), .C(n5717), .D(n1), 
         .Z(n8845)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4521_4_lut.init = 16'hc0ca;
    LUT4 i4523_4_lut (.A(n3930[11]), .B(quad_set[11]), .C(n5717), .D(n1), 
         .Z(n8847)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4523_4_lut.init = 16'hc0ca;
    LUT4 i4525_4_lut (.A(n3930[10]), .B(quad_set[10]), .C(n5717), .D(n1), 
         .Z(n8849)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4525_4_lut.init = 16'hc0ca;
    LUT4 i4527_4_lut (.A(n3930[9]), .B(quad_set[9]), .C(n5717), .D(n1), 
         .Z(n8851)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4527_4_lut.init = 16'hc0ca;
    LUT4 i4529_4_lut (.A(n3930[8]), .B(quad_set[8]), .C(n5717), .D(n1), 
         .Z(n8853)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4529_4_lut.init = 16'hc0ca;
    LUT4 i4531_4_lut (.A(n3930[7]), .B(quad_set[7]), .C(n5717), .D(n1), 
         .Z(n8855)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4531_4_lut.init = 16'hc0ca;
    LUT4 i4533_4_lut (.A(n3930[6]), .B(quad_set[6]), .C(n5717), .D(n1), 
         .Z(n8857)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4533_4_lut.init = 16'hc0ca;
    LUT4 i4535_4_lut (.A(n3930[5]), .B(quad_set[5]), .C(n5717), .D(n1), 
         .Z(n8859)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4535_4_lut.init = 16'hc0ca;
    LUT4 i4537_4_lut (.A(n3930[4]), .B(quad_set[4]), .C(n5717), .D(n1), 
         .Z(n8861)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4537_4_lut.init = 16'hc0ca;
    LUT4 i4539_4_lut (.A(n3930[3]), .B(quad_set[3]), .C(n5717), .D(n1), 
         .Z(n8863)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4539_4_lut.init = 16'hc0ca;
    LUT4 i4541_4_lut (.A(n3930[2]), .B(quad_set[2]), .C(n5717), .D(n1), 
         .Z(n8865)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4541_4_lut.init = 16'hc0ca;
    LUT4 i4543_4_lut (.A(n3930[1]), .B(quad_set[1]), .C(n5717), .D(n1), 
         .Z(n8867)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4543_4_lut.init = 16'hc0ca;
    
endmodule
//
// Verilog Description of module \servo(UART_ADDRESS_WIDTH=4) 
//

module \servo(UART_ADDRESS_WIDTH=4)  (pin_io_out_2, pin_io_out_1, n30043, 
            mode, \pin_intrpt[0] , clk, clk_enable_232, n30185, \spi_data_r[0] , 
            Phase_r, clk_enable_234, pin_io_out_9, \quad_b[0] , mode_adj_655, 
            \spi_cmd_r[2] , \spi_cmd_r[0] , n23732, pin_io_out_8, \quad_a[0] , 
            \uart_slot_en[3] , \uart_slot_en[0] , n8, pin_io_out_3, 
            \pin_intrpt[1] ) /* synthesis syn_module_defined=1 */ ;
    input pin_io_out_2;
    input pin_io_out_1;
    input n30043;
    output mode;
    output \pin_intrpt[0] ;
    input clk;
    input clk_enable_232;
    input n30185;
    input \spi_data_r[0] ;
    output Phase_r;
    input clk_enable_234;
    input pin_io_out_9;
    output \quad_b[0] ;
    input [2:0]mode_adj_655;
    input \spi_cmd_r[2] ;
    input \spi_cmd_r[0] ;
    output n23732;
    input pin_io_out_8;
    output \quad_a[0] ;
    input \uart_slot_en[3] ;
    input \uart_slot_en[0] ;
    output n8;
    input pin_io_out_3;
    output \pin_intrpt[1] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    
    wire n7212;
    
    LUT4 Select_2918_i3_4_lut (.A(pin_io_out_2), .B(pin_io_out_1), .C(n30043), 
         .D(mode), .Z(\pin_intrpt[0] )) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam Select_2918_i3_4_lut.init = 16'heca0;
    FD1P3IX mode_76 (.D(\spi_data_r[0] ), .SP(clk_enable_232), .CD(n30185), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=408, LSE_RLINE=443 */ ;   // c:/s_links/sources/slot_cards/servo.v(66[8] 74[4])
    defparam mode_76.GSR = "DISABLED";
    FD1P3IX Phase_r_77 (.D(\spi_data_r[0] ), .SP(clk_enable_234), .CD(n30185), 
            .CK(clk), .Q(Phase_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=408, LSE_RLINE=443 */ ;   // c:/s_links/sources/slot_cards/servo.v(77[8] 85[4])
    defparam Phase_r_77.GSR = "DISABLED";
    LUT4 i3000_2_lut (.A(pin_io_out_9), .B(n7212), .Z(\quad_b[0] )) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/servo.v(56[8:18])
    defparam i3000_2_lut.init = 16'h8888;
    LUT4 i2916_4_lut (.A(mode_adj_655[1]), .B(mode), .C(mode_adj_655[0]), 
         .D(mode_adj_655[2]), .Z(n7212)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/s_links/sources/slot_cards/servo.v(55[8:18])
    defparam i2916_4_lut.init = 16'hccdc;
    LUT4 i19108_2_lut (.A(\spi_cmd_r[2] ), .B(\spi_cmd_r[0] ), .Z(n23732)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i19108_2_lut.init = 16'heeee;
    LUT4 i2999_2_lut (.A(pin_io_out_8), .B(n7212), .Z(\quad_a[0] )) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/servo.v(55[8:18])
    defparam i2999_2_lut.init = 16'h8888;
    LUT4 i3_3_lut (.A(\uart_slot_en[3] ), .B(\uart_slot_en[0] ), .C(mode), 
         .Z(n8)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i3_3_lut.init = 16'h4040;
    LUT4 Select_2917_i3_4_lut (.A(pin_io_out_3), .B(pin_io_out_2), .C(n30043), 
         .D(mode), .Z(\pin_intrpt[1] )) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam Select_2917_i3_4_lut.init = 16'heca0;
    
endmodule
//
// Verilog Description of module \otm_dac(DEV_ID=3) 
//

module \otm_dac(DEV_ID=3)  (clk, clk_enable_255, n30185, \spi_data_r[0] , 
            mode, clk_enable_260, NSL, n30082, n7167) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input clk_enable_255;
    input n30185;
    input \spi_data_r[0] ;
    output mode;
    input clk_enable_260;
    input NSL;
    input n30082;
    output n7167;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    
    wire LASER_CNTRL_r;
    
    FD1P3IX LASER_CNTRL_r_31 (.D(\spi_data_r[0] ), .SP(clk_enable_255), 
            .CD(n30185), .CK(clk), .Q(LASER_CNTRL_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=566, LSE_RLINE=584 */ ;   // c:/s_links/sources/otm_dac.v(47[8] 55[4])
    defparam LASER_CNTRL_r_31.GSR = "DISABLED";
    FD1P3IX mode_30 (.D(\spi_data_r[0] ), .SP(clk_enable_260), .CD(n30185), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=566, LSE_RLINE=584 */ ;   // c:/s_links/sources/otm_dac.v(36[8] 44[4])
    defparam mode_30.GSR = "DISABLED";
    LUT4 Select_2829_i3_4_lut (.A(NSL), .B(LASER_CNTRL_r), .C(n30082), 
         .D(mode), .Z(n7167)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;
    defparam Select_2829_i3_4_lut.init = 16'hce0a;
    
endmodule
//
// Verilog Description of module \stepper(DEV_ID=5,UART_ADDRESS_WIDTH=4) 
//

module \stepper(DEV_ID=5,UART_ADDRESS_WIDTH=4)  (clk_1MHz, n30185, clk, 
            reset_r, clk_enable_38, n29994, clk_enable_627, \spi_data_r[0] , 
            GND_net, pin_io_c_58, n30149, spi_data_out_r_39__N_5540, 
            resetn_c, digital_output_r, clk_enable_242, n28551, spi_data_out_r_39__N_5580, 
            spi_data_out_r_39__N_5877, \spi_data_r[1] , \spi_data_r[2] , 
            n47, NSL, \uart_slot_en[2] , \uart_slot_en[3] , n10696, 
            \quad_homing[0] , pin_io_c_54, n25885, pin_io_out_59, \quad_b[5] , 
            UC_TXD0_c, OW_ID_N_5833, OW_ID_N_5839, n30049, \uart_slot_en[0] , 
            \quad_a[5] , n30047, n30087, \pin_intrpt[17] , n7262, 
            pin_io_c_52, \pin_intrpt[15] , pin_io_c_53, \pin_intrpt[16] , 
            ENC_O_N_5841) /* synthesis syn_module_defined=1 */ ;
    input clk_1MHz;
    input n30185;
    input clk;
    output reset_r;
    input clk_enable_38;
    input n29994;
    input clk_enable_627;
    input \spi_data_r[0] ;
    input GND_net;
    input pin_io_c_58;
    output n30149;
    output [39:0]spi_data_out_r_39__N_5540;
    input resetn_c;
    output digital_output_r;
    input clk_enable_242;
    input n28551;
    output spi_data_out_r_39__N_5580;
    input spi_data_out_r_39__N_5877;
    input \spi_data_r[1] ;
    input \spi_data_r[2] ;
    input n47;
    output NSL;
    input \uart_slot_en[2] ;
    input \uart_slot_en[3] ;
    output n10696;
    input \quad_homing[0] ;
    input pin_io_c_54;
    output n25885;
    input pin_io_out_59;
    output \quad_b[5] ;
    input UC_TXD0_c;
    output OW_ID_N_5833;
    output OW_ID_N_5839;
    input n30049;
    input \uart_slot_en[0] ;
    output \quad_a[5] ;
    output n30047;
    output n30087;
    output \pin_intrpt[17] ;
    output n7262;
    input pin_io_c_52;
    output \pin_intrpt[15] ;
    input pin_io_c_53;
    output \pin_intrpt[16] ;
    output ENC_O_N_5841;
    
    wire clk_1MHz /* synthesis SET_AS_NETWORK=clk_1MHz, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(136[6:14])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire \pin_intrpt[17]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[17] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    
    wire MA_Temp, clk_1MHz_enable_3, MA_Temp_N_5859;
    wire [51:0]SLO_buf;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire SLO_buf_51__N_5730;
    wire [51:0]SLO;   // c:/s_links/sources/slot_cards/stepper.v(63[12:15])
    wire [7:0]Cnt;   // c:/s_links/sources/slot_cards/stepper.v(62[11:14])
    
    wire clk_1MHz_enable_34;
    wire [7:0]n199;
    wire [2:0]mode;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    wire clk_enable_1057, prev_MA_Temp, prev_MA;
    wire [39:0]spi_data_out_r_39__N_5791;
    wire [11:0]n93;
    wire [11:0]n53;
    
    wire n30111, n26369, n30067, n30133, n30132, n18602, clk_1MHz_enable_69, 
        n12542, n18532;
    wire [31:0]n153;
    
    wire n4, n28591, n28592;
    wire [11:0]Cnt_NSL;   // c:/s_links/sources/slot_cards/stepper.v(61[12:19])
    
    wire n28320, n30066, n30057, n30006, NSL_N_5872, n21963, n21962, 
        n21961, n21960, n22019, n22018, n22017, n22016, n22015, 
        n22014, n30115, n25174, n30112, n18446, n26309, OW_ID_N_5834, 
        n28368, n30191, n30116;
    
    FD1P3IX MA_Temp_483 (.D(MA_Temp_N_5859), .SP(clk_1MHz_enable_3), .CD(n30185), 
            .CK(clk_1MHz), .Q(MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam MA_Temp_483.GSR = "DISABLED";
    FD1P3AX SLO_buf__i1 (.D(SLO[0]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i1.GSR = "DISABLED";
    FD1P3IX Cnt__i0 (.D(n199[0]), .SP(clk_1MHz_enable_34), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i0.GSR = "DISABLED";
    FD1P3IX reset_r_491 (.D(n29994), .SP(clk_enable_38), .CD(n30185), 
            .CK(clk), .Q(reset_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam reset_r_491.GSR = "DISABLED";
    FD1P3IX mode__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_627), .CD(n30185), 
            .CK(clk), .Q(mode[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i0.GSR = "DISABLED";
    FD1P3IX SLO__i1 (.D(pin_io_c_58), .SP(clk_enable_1057), .CD(GND_net), 
            .CK(clk), .Q(SLO[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i1.GSR = "DISABLED";
    FD1S3AX prev_MA_Temp_487 (.D(MA_Temp), .CK(clk), .Q(prev_MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam prev_MA_Temp_487.GSR = "DISABLED";
    FD1S3AX prev_MA_489 (.D(n30149), .CK(clk), .Q(prev_MA)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam prev_MA_489.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i0 (.D(spi_data_out_r_39__N_5791[0]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i0.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1783__i0 (.D(n53[0]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783__i0.GSR = "DISABLED";
    LUT4 i24147_4_lut_4_lut (.A(mode[2]), .B(n30111), .C(n26369), .D(n30067), 
         .Z(clk_enable_1057)) /* synthesis lut_function=(!(A (B+(D))+!A ((D)+!C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i24147_4_lut_4_lut.init = 16'h0072;
    FD1P3IX digital_output_r_492 (.D(n28551), .SP(clk_enable_242), .CD(n30185), 
            .CK(clk), .Q(digital_output_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam digital_output_r_492.GSR = "DISABLED";
    FD1S3IX i168_494 (.D(spi_data_out_r_39__N_5877), .CK(clk), .CD(n30185), 
            .Q(spi_data_out_r_39__N_5580)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam i168_494.GSR = "DISABLED";
    LUT4 i14069_3_lut_4_lut (.A(n30133), .B(n30132), .C(resetn_c), .D(n18602), 
         .Z(clk_1MHz_enable_69)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i14069_3_lut_4_lut.init = 16'h70f0;
    LUT4 i24106_2_lut_3_lut_4_lut (.A(prev_MA), .B(n30149), .C(n30111), 
         .D(mode[2]), .Z(n12542)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i24106_2_lut_3_lut_4_lut.init = 16'h0400;
    LUT4 i13007_2_lut_3_lut (.A(n18532), .B(n18602), .C(n153[0]), .Z(n199[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13007_2_lut_3_lut.init = 16'h7070;
    FD1P3IX Cnt__i7 (.D(n199[7]), .SP(clk_1MHz_enable_34), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i7.GSR = "DISABLED";
    LUT4 i13549_2_lut_3_lut (.A(n18532), .B(n18602), .C(n153[7]), .Z(n199[7])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13549_2_lut_3_lut.init = 16'h7070;
    FD1P3IX Cnt__i6 (.D(n199[6]), .SP(clk_1MHz_enable_34), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i6.GSR = "DISABLED";
    FD1P3IX Cnt__i5 (.D(n199[5]), .SP(clk_1MHz_enable_34), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i5.GSR = "DISABLED";
    FD1P3IX Cnt__i4 (.D(n199[4]), .SP(clk_1MHz_enable_34), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i4.GSR = "DISABLED";
    LUT4 i13548_2_lut_3_lut (.A(n18532), .B(n18602), .C(n153[6]), .Z(n199[6])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13548_2_lut_3_lut.init = 16'h7070;
    FD1P3IX Cnt__i3 (.D(n199[3]), .SP(clk_1MHz_enable_34), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i3.GSR = "DISABLED";
    FD1P3IX Cnt__i2 (.D(n199[2]), .SP(clk_1MHz_enable_34), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i1 (.D(n199[1]), .SP(clk_1MHz_enable_34), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i1.GSR = "DISABLED";
    FD1P3AX SLO_buf__i46 (.D(SLO[45]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i46.GSR = "DISABLED";
    FD1P3AX SLO_buf__i45 (.D(SLO[44]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i45.GSR = "DISABLED";
    FD1P3AX SLO_buf__i44 (.D(SLO[43]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i44.GSR = "DISABLED";
    FD1P3AX SLO_buf__i43 (.D(SLO[42]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i43.GSR = "DISABLED";
    FD1P3AX SLO_buf__i42 (.D(SLO[41]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i42.GSR = "DISABLED";
    FD1P3AX SLO_buf__i41 (.D(SLO[40]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i41.GSR = "DISABLED";
    FD1P3AX SLO_buf__i40 (.D(SLO[39]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i40.GSR = "DISABLED";
    FD1P3AX SLO_buf__i39 (.D(SLO[38]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i39.GSR = "DISABLED";
    FD1P3AX SLO_buf__i38 (.D(SLO[37]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i38.GSR = "DISABLED";
    FD1P3AX SLO_buf__i37 (.D(SLO[36]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i37.GSR = "DISABLED";
    FD1P3AX SLO_buf__i36 (.D(SLO[35]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i36.GSR = "DISABLED";
    FD1P3AX SLO_buf__i35 (.D(SLO[34]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i35.GSR = "DISABLED";
    FD1P3AX SLO_buf__i34 (.D(SLO[33]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i34.GSR = "DISABLED";
    FD1P3AX SLO_buf__i33 (.D(SLO[32]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i33.GSR = "DISABLED";
    FD1P3AX SLO_buf__i32 (.D(SLO[31]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i32.GSR = "DISABLED";
    FD1P3AX SLO_buf__i31 (.D(SLO[30]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i31.GSR = "DISABLED";
    FD1P3AX SLO_buf__i30 (.D(SLO[29]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i30.GSR = "DISABLED";
    FD1P3AX SLO_buf__i29 (.D(SLO[28]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i29.GSR = "DISABLED";
    FD1P3AX SLO_buf__i28 (.D(SLO[27]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i28.GSR = "DISABLED";
    FD1P3AX SLO_buf__i27 (.D(SLO[26]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i27.GSR = "DISABLED";
    FD1P3AX SLO_buf__i26 (.D(SLO[25]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i26.GSR = "DISABLED";
    FD1P3AX SLO_buf__i25 (.D(SLO[24]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i25.GSR = "DISABLED";
    FD1P3AX SLO_buf__i24 (.D(SLO[23]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i24.GSR = "DISABLED";
    FD1P3AX SLO_buf__i23 (.D(SLO[22]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i23.GSR = "DISABLED";
    FD1P3AX SLO_buf__i22 (.D(SLO[21]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i22.GSR = "DISABLED";
    FD1P3AX SLO_buf__i21 (.D(SLO[20]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i21.GSR = "DISABLED";
    FD1P3AX SLO_buf__i20 (.D(SLO[19]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i20.GSR = "DISABLED";
    FD1P3AX SLO_buf__i19 (.D(SLO[18]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i19.GSR = "DISABLED";
    FD1P3AX SLO_buf__i18 (.D(SLO[17]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i18.GSR = "DISABLED";
    FD1P3AX SLO_buf__i17 (.D(SLO[16]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i17.GSR = "DISABLED";
    FD1P3AX SLO_buf__i16 (.D(SLO[15]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i16.GSR = "DISABLED";
    FD1P3AX SLO_buf__i15 (.D(SLO[14]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i15.GSR = "DISABLED";
    FD1P3AX SLO_buf__i14 (.D(SLO[13]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i14.GSR = "DISABLED";
    FD1P3AX SLO_buf__i13 (.D(SLO[12]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i13.GSR = "DISABLED";
    FD1P3AX SLO_buf__i12 (.D(SLO[11]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i12.GSR = "DISABLED";
    FD1P3AX SLO_buf__i11 (.D(SLO[10]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i11.GSR = "DISABLED";
    FD1P3AX SLO_buf__i10 (.D(SLO[9]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i10.GSR = "DISABLED";
    FD1P3AX SLO_buf__i9 (.D(SLO[8]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i9.GSR = "DISABLED";
    FD1P3AX SLO_buf__i8 (.D(SLO[7]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i8.GSR = "DISABLED";
    FD1P3AX SLO_buf__i7 (.D(SLO[6]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i7.GSR = "DISABLED";
    FD1P3AX SLO_buf__i6 (.D(SLO[5]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i6.GSR = "DISABLED";
    FD1P3AX SLO_buf__i5 (.D(SLO[4]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i5.GSR = "DISABLED";
    FD1P3AX SLO_buf__i4 (.D(SLO[3]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i4.GSR = "DISABLED";
    FD1P3AX SLO_buf__i3 (.D(SLO[2]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i3.GSR = "DISABLED";
    FD1P3AX SLO_buf__i2 (.D(SLO[1]), .SP(SLO_buf_51__N_5730), .CK(clk), 
            .Q(SLO_buf[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i2.GSR = "DISABLED";
    LUT4 SLO_buf_51__I_214_2_lut (.A(prev_MA_Temp), .B(MA_Temp), .Z(SLO_buf_51__N_5730)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[5:38])
    defparam SLO_buf_51__I_214_2_lut.init = 16'h2222;
    LUT4 i1_4_lut (.A(mode[1]), .B(mode[0]), .C(Cnt[4]), .D(n4), .Z(n26369)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut.init = 16'h8880;
    LUT4 i13547_2_lut_3_lut (.A(n18532), .B(n18602), .C(n153[5]), .Z(n199[5])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13547_2_lut_3_lut.init = 16'h7070;
    LUT4 i13546_2_lut_3_lut (.A(n18532), .B(n18602), .C(n153[4]), .Z(n199[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13546_2_lut_3_lut.init = 16'h7070;
    FD1P3IX mode__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_627), .CD(n30185), 
            .CK(clk), .Q(mode[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i1.GSR = "DISABLED";
    FD1P3IX mode__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_627), .CD(n30185), 
            .CK(clk), .Q(mode[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i2.GSR = "DISABLED";
    PFUMX MA_Temp_I_229 (.BLUT(n28591), .ALUT(n28592), .C0(n18602), .Z(MA_Temp_N_5859)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;
    LUT4 i13545_2_lut_3_lut (.A(n18532), .B(n18602), .C(n153[3]), .Z(n199[3])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13545_2_lut_3_lut.init = 16'h7070;
    LUT4 i13544_2_lut_3_lut (.A(n18532), .B(n18602), .C(n153[2]), .Z(n199[2])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13544_2_lut_3_lut.init = 16'h7070;
    FD1S3AX spi_data_out_r_i1 (.D(spi_data_out_r_39__N_5791[1]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(spi_data_out_r_39__N_5791[2]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(spi_data_out_r_39__N_5791[3]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(spi_data_out_r_39__N_5791[4]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(spi_data_out_r_39__N_5791[5]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(spi_data_out_r_39__N_5791[6]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(spi_data_out_r_39__N_5791[7]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(spi_data_out_r_39__N_5791[8]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(spi_data_out_r_39__N_5791[9]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(spi_data_out_r_39__N_5791[10]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(spi_data_out_r_39__N_5791[11]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(spi_data_out_r_39__N_5791[12]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(spi_data_out_r_39__N_5791[13]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(spi_data_out_r_39__N_5791[14]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(spi_data_out_r_39__N_5791[15]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i16 (.D(SLO_buf[30]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i17 (.D(SLO_buf[31]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i18 (.D(SLO_buf[32]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i19 (.D(SLO_buf[33]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i20 (.D(SLO_buf[34]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i21 (.D(SLO_buf[35]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i22 (.D(SLO_buf[36]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i23 (.D(SLO_buf[37]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i24 (.D(SLO_buf[38]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i25 (.D(SLO_buf[39]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i26 (.D(SLO_buf[40]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i27 (.D(SLO_buf[41]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i28 (.D(SLO_buf[42]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i29 (.D(SLO_buf[43]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i30 (.D(SLO_buf[44]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i31 (.D(SLO_buf[45]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(spi_data_out_r_39__N_5791[32]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i33 (.D(spi_data_out_r_39__N_5791[33]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i33.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i34 (.D(spi_data_out_r_39__N_5791[34]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i34.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i35 (.D(spi_data_out_r_39__N_5791[35]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5540[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i35.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i36 (.D(SLO_buf[10]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i36.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i37 (.D(SLO_buf[11]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i37.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i38 (.D(SLO_buf[12]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i38.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i39 (.D(SLO_buf[13]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5540[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i39.GSR = "DISABLED";
    LUT4 i13543_2_lut_3_lut (.A(n18532), .B(n18602), .C(n153[1]), .Z(n199[1])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13543_2_lut_3_lut.init = 16'h7070;
    FD1P3AX Cnt_NSL_1783__i1 (.D(n53[1]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783__i1.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1783__i2 (.D(n53[2]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783__i2.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1783__i3 (.D(n53[3]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783__i3.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1783__i4 (.D(n53[4]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783__i4.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1783__i5 (.D(n53[5]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783__i5.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1783__i6 (.D(n53[6]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783__i6.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1783__i7 (.D(n53[7]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783__i7.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1783__i8 (.D(n53[8]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783__i8.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1783__i9 (.D(n53[9]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783__i9.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1783__i10 (.D(n53[10]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783__i10.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1783__i11 (.D(n53[11]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783__i11.GSR = "DISABLED";
    LUT4 mux_158_i1_3_lut (.A(SLO_buf[14]), .B(SLO_buf[4]), .C(n47), .Z(spi_data_out_r_39__N_5791[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i1_3_lut.init = 16'hcaca;
    LUT4 i23901_1_lut_4_lut (.A(MA_Temp), .B(n18532), .C(n28320), .D(n30066), 
         .Z(n28592)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A (B+((D)+!C)))) */ ;
    defparam i23901_1_lut_4_lut.init = 16'h2212;
    LUT4 i23992_4_lut (.A(NSL), .B(n30057), .C(n18602), .D(n30006), 
         .Z(NSL_N_5872)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C+(D))))) */ ;
    defparam i23992_4_lut.init = 16'h3b37;
    CCU2D add_564_9 (.A0(Cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21963), 
          .S0(n153[7]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_9.INIT0 = 16'h5aaa;
    defparam add_564_9.INIT1 = 16'h0000;
    defparam add_564_9.INJECT1_0 = "NO";
    defparam add_564_9.INJECT1_1 = "NO";
    CCU2D add_564_7 (.A0(Cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21962), 
          .COUT(n21963), .S0(n153[5]), .S1(n153[6]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_7.INIT0 = 16'h5aaa;
    defparam add_564_7.INIT1 = 16'h5aaa;
    defparam add_564_7.INJECT1_0 = "NO";
    defparam add_564_7.INJECT1_1 = "NO";
    CCU2D add_564_5 (.A0(Cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21961), 
          .COUT(n21962), .S0(n153[3]), .S1(n153[4]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_5.INIT0 = 16'h5aaa;
    defparam add_564_5.INIT1 = 16'h5aaa;
    defparam add_564_5.INJECT1_0 = "NO";
    defparam add_564_5.INJECT1_1 = "NO";
    CCU2D add_564_3 (.A0(Cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21960), 
          .COUT(n21961), .S0(n153[1]), .S1(n153[2]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_3.INIT0 = 16'h5aaa;
    defparam add_564_3.INIT1 = 16'h5aaa;
    defparam add_564_3.INJECT1_0 = "NO";
    defparam add_564_3.INJECT1_1 = "NO";
    CCU2D add_564_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n21960), 
          .S1(n153[0]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_1.INIT0 = 16'hF000;
    defparam add_564_1.INIT1 = 16'h5555;
    defparam add_564_1.INJECT1_0 = "NO";
    defparam add_564_1.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1783_add_4_13 (.A0(Cnt_NSL[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n22019), .S0(n53[11]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783_add_4_13.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1783_add_4_13.INIT1 = 16'h0000;
    defparam Cnt_NSL_1783_add_4_13.INJECT1_0 = "NO";
    defparam Cnt_NSL_1783_add_4_13.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1783_add_4_11 (.A0(Cnt_NSL[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Cnt_NSL[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22018), .COUT(n22019), .S0(n53[9]), .S1(n53[10]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783_add_4_11.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1783_add_4_11.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1783_add_4_11.INJECT1_0 = "NO";
    defparam Cnt_NSL_1783_add_4_11.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1783_add_4_9 (.A0(Cnt_NSL[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Cnt_NSL[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22017), .COUT(n22018), .S0(n53[7]), .S1(n53[8]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783_add_4_9.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1783_add_4_9.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1783_add_4_9.INJECT1_0 = "NO";
    defparam Cnt_NSL_1783_add_4_9.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1783_add_4_7 (.A0(n93[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n22016), .COUT(n22017), .S0(n53[5]), .S1(n53[6]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783_add_4_7.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1783_add_4_7.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1783_add_4_7.INJECT1_0 = "NO";
    defparam Cnt_NSL_1783_add_4_7.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1783_add_4_5 (.A0(n93[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n22015), .COUT(n22016), .S0(n53[3]), .S1(n53[4]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783_add_4_5.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1783_add_4_5.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1783_add_4_5.INJECT1_0 = "NO";
    defparam Cnt_NSL_1783_add_4_5.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1783_add_4_3 (.A0(n93[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n22014), .COUT(n22015), .S0(n53[1]), .S1(n53[2]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783_add_4_3.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1783_add_4_3.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1783_add_4_3.INJECT1_0 = "NO";
    defparam Cnt_NSL_1783_add_4_3.INJECT1_1 = "NO";
    LUT4 i12758_2_lut (.A(\uart_slot_en[2] ), .B(\uart_slot_en[3] ), .Z(n10696)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12758_2_lut.init = 16'h8888;
    CCU2D Cnt_NSL_1783_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n30132), .B1(n30133), .C1(n93[0]), .D1(GND_net), 
          .COUT(n22014), .S1(n53[0]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1783_add_4_1.INIT0 = 16'hF000;
    defparam Cnt_NSL_1783_add_4_1.INIT1 = 16'h8787;
    defparam Cnt_NSL_1783_add_4_1.INJECT1_0 = "NO";
    defparam Cnt_NSL_1783_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(\quad_homing[0] ), .B(pin_io_c_54), .Z(n25885)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(74[8:17])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_847 (.A(n30115), .B(n25174), .C(n30112), .D(mode[2]), 
         .Z(n18532)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(107[27:54])
    defparam i1_4_lut_adj_847.init = 16'hffef;
    LUT4 i1_3_lut (.A(Cnt[5]), .B(n18446), .C(Cnt[4]), .Z(n25174)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_adj_848 (.A(n30115), .B(n18446), .C(n26309), .D(Cnt[4]), 
         .Z(n18602)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_848.init = 16'hfefa;
    LUT4 mux_158_i2_3_lut (.A(SLO_buf[15]), .B(SLO_buf[5]), .C(n47), .Z(spi_data_out_r_39__N_5791[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i2_3_lut.init = 16'hcaca;
    LUT4 mux_158_i3_3_lut (.A(SLO_buf[16]), .B(SLO_buf[6]), .C(n47), .Z(spi_data_out_r_39__N_5791[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i3_3_lut.init = 16'hcaca;
    LUT4 mux_158_i4_3_lut (.A(SLO_buf[17]), .B(SLO_buf[7]), .C(n47), .Z(spi_data_out_r_39__N_5791[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i4_3_lut.init = 16'hcaca;
    LUT4 mux_158_i5_3_lut (.A(SLO_buf[18]), .B(SLO_buf[8]), .C(n47), .Z(spi_data_out_r_39__N_5791[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i5_3_lut.init = 16'hcaca;
    LUT4 mux_158_i6_3_lut (.A(SLO_buf[19]), .B(SLO_buf[9]), .C(n47), .Z(spi_data_out_r_39__N_5791[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i6_3_lut.init = 16'hcaca;
    LUT4 mux_158_i7_3_lut (.A(SLO_buf[20]), .B(SLO_buf[10]), .C(n47), 
         .Z(spi_data_out_r_39__N_5791[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i7_3_lut.init = 16'hcaca;
    LUT4 mux_158_i8_3_lut (.A(SLO_buf[21]), .B(SLO_buf[11]), .C(n47), 
         .Z(spi_data_out_r_39__N_5791[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i8_3_lut.init = 16'hcaca;
    LUT4 mux_158_i9_3_lut (.A(SLO_buf[22]), .B(SLO_buf[12]), .C(n47), 
         .Z(spi_data_out_r_39__N_5791[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i9_3_lut.init = 16'hcaca;
    LUT4 mux_158_i10_3_lut (.A(SLO_buf[23]), .B(SLO_buf[13]), .C(n47), 
         .Z(spi_data_out_r_39__N_5791[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i10_3_lut.init = 16'hcaca;
    LUT4 mux_158_i11_3_lut (.A(SLO_buf[24]), .B(SLO_buf[14]), .C(n47), 
         .Z(spi_data_out_r_39__N_5791[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i11_3_lut.init = 16'hcaca;
    LUT4 mux_158_i12_3_lut (.A(SLO_buf[25]), .B(SLO_buf[15]), .C(n47), 
         .Z(spi_data_out_r_39__N_5791[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i12_3_lut.init = 16'hcaca;
    LUT4 mux_158_i13_3_lut (.A(SLO_buf[26]), .B(SLO_buf[16]), .C(n47), 
         .Z(spi_data_out_r_39__N_5791[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i13_3_lut.init = 16'hcaca;
    LUT4 mux_158_i14_3_lut (.A(SLO_buf[27]), .B(SLO_buf[17]), .C(n47), 
         .Z(spi_data_out_r_39__N_5791[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i14_3_lut.init = 16'hcaca;
    LUT4 mux_158_i15_3_lut (.A(SLO_buf[28]), .B(SLO_buf[18]), .C(n47), 
         .Z(spi_data_out_r_39__N_5791[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i15_3_lut.init = 16'hcaca;
    LUT4 mux_158_i16_3_lut (.A(SLO_buf[29]), .B(SLO_buf[19]), .C(n47), 
         .Z(spi_data_out_r_39__N_5791[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i16_3_lut.init = 16'hcaca;
    LUT4 mux_158_i33_3_lut (.A(SLO_buf[6]), .B(SLO_buf[0]), .C(n47), .Z(spi_data_out_r_39__N_5791[32])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i33_3_lut.init = 16'hcaca;
    LUT4 i2993_2_lut_4_lut (.A(mode[2]), .B(mode[0]), .C(mode[1]), .D(pin_io_out_59), 
         .Z(\quad_b[5] )) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i2993_2_lut_4_lut.init = 16'h0400;
    LUT4 mux_158_i34_3_lut (.A(SLO_buf[7]), .B(SLO_buf[1]), .C(n47), .Z(spi_data_out_r_39__N_5791[33])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i34_3_lut.init = 16'hcaca;
    LUT4 mux_158_i35_3_lut (.A(SLO_buf[8]), .B(SLO_buf[2]), .C(n47), .Z(spi_data_out_r_39__N_5791[34])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i35_3_lut.init = 16'hcaca;
    LUT4 digital_output_r_I_0_547_3_lut (.A(digital_output_r), .B(UC_TXD0_c), 
         .C(OW_ID_N_5834), .Z(OW_ID_N_5833)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[16] 91[59])
    defparam digital_output_r_I_0_547_3_lut.init = 16'hcaca;
    LUT4 mux_158_i36_3_lut (.A(SLO_buf[9]), .B(SLO_buf[3]), .C(n47), .Z(spi_data_out_r_39__N_5791[35])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i36_3_lut.init = 16'hcaca;
    LUT4 i24088_4_lut (.A(OW_ID_N_5834), .B(mode[1]), .C(mode[0]), .D(mode[2]), 
         .Z(OW_ID_N_5839)) /* synthesis lut_function=(!(A+!((C+(D))+!B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[8:13])
    defparam i24088_4_lut.init = 16'h5551;
    LUT4 i4_4_lut (.A(mode[0]), .B(mode[2]), .C(n30049), .D(n28368), 
         .Z(OW_ID_N_5834)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i4_4_lut.init = 16'h0020;
    LUT4 i23666_2_lut (.A(\uart_slot_en[0] ), .B(mode[1]), .Z(n28368)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23666_2_lut.init = 16'heeee;
    LUT4 i2992_2_lut_4_lut (.A(mode[2]), .B(mode[0]), .C(mode[1]), .D(pin_io_c_58), 
         .Z(\quad_a[5] )) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i2992_2_lut_4_lut.init = 16'h0400;
    LUT4 i13240_2_lut_rep_791 (.A(Cnt[4]), .B(Cnt[1]), .Z(n30191)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13240_2_lut_rep_791.init = 16'h8888;
    LUT4 i23618_2_lut_3_lut (.A(Cnt[4]), .B(Cnt[1]), .C(Cnt[5]), .Z(n28320)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i23618_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_606_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(n30066), 
         .D(Cnt[5]), .Z(n30006)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_rep_606_3_lut_4_lut.init = 16'hfff7;
    LUT4 i24103_2_lut_3_lut_4_lut (.A(n30057), .B(resetn_c), .C(n18602), 
         .D(n18532), .Z(clk_1MHz_enable_3)) /* synthesis lut_function=(!(A (C (D))+!A (B+(C (D))))) */ ;
    defparam i24103_2_lut_3_lut_4_lut.init = 16'h0bbb;
    LUT4 i1_2_lut_3_lut (.A(Cnt[5]), .B(n30066), .C(Cnt[1]), .Z(n4)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(133[16:19])
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i23900_1_lut_2_lut_3_lut_4_lut (.A(Cnt[5]), .B(n30066), .C(MA_Temp), 
         .D(n30191), .Z(n28591)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(133[16:19])
    defparam i23900_1_lut_2_lut_3_lut_4_lut.init = 16'he1f0;
    FD1P3IX SLO__i45 (.D(SLO[43]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i45.GSR = "DISABLED";
    FD1P3IX SLO__i46 (.D(SLO[44]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i46.GSR = "DISABLED";
    FD1P3IX SLO__i43 (.D(SLO[41]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i43.GSR = "DISABLED";
    FD1P3IX SLO__i44 (.D(SLO[42]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i44.GSR = "DISABLED";
    FD1P3IX SLO__i33 (.D(SLO[31]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i33.GSR = "DISABLED";
    FD1P3IX SLO__i37 (.D(SLO[35]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i37.GSR = "DISABLED";
    FD1P3IX SLO__i40 (.D(SLO[38]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i40.GSR = "DISABLED";
    FD1P3IX SLO__i34 (.D(SLO[32]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i34.GSR = "DISABLED";
    FD1P3IX SLO__i38 (.D(SLO[36]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i38.GSR = "DISABLED";
    FD1P3IX SLO__i41 (.D(SLO[39]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i41.GSR = "DISABLED";
    FD1P3IX SLO__i31 (.D(SLO[29]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i31.GSR = "DISABLED";
    FD1P3IX SLO__i35 (.D(SLO[33]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i35.GSR = "DISABLED";
    FD1P3IX SLO__i32 (.D(SLO[30]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i32.GSR = "DISABLED";
    FD1P3IX SLO__i36 (.D(SLO[34]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i36.GSR = "DISABLED";
    FD1P3IX SLO__i39 (.D(SLO[37]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i39.GSR = "DISABLED";
    FD1P3IX SLO__i42 (.D(SLO[40]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i42.GSR = "DISABLED";
    FD1P3IX SLO__i21 (.D(SLO[19]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i21.GSR = "DISABLED";
    FD1P3IX SLO__i25 (.D(SLO[23]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i25.GSR = "DISABLED";
    FD1P3IX SLO__i28 (.D(SLO[26]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i28.GSR = "DISABLED";
    FD1P3IX SLO__i22 (.D(SLO[20]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i22.GSR = "DISABLED";
    FD1P3IX SLO__i26 (.D(SLO[24]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i26.GSR = "DISABLED";
    FD1P3IX SLO__i29 (.D(SLO[27]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i29.GSR = "DISABLED";
    FD1P3IX SLO__i20 (.D(SLO[18]), .SP(clk_enable_1057), .CD(GND_net), 
            .CK(clk), .Q(SLO[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i20.GSR = "DISABLED";
    FD1P3IX SLO__i23 (.D(SLO[21]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i23.GSR = "DISABLED";
    FD1P3IX SLO__i24 (.D(SLO[22]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i24.GSR = "DISABLED";
    FD1P3IX SLO__i27 (.D(SLO[25]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i27.GSR = "DISABLED";
    FD1P3IX SLO__i30 (.D(SLO[28]), .SP(clk_enable_1057), .CD(n12542), 
            .CK(clk), .Q(SLO[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i30.GSR = "DISABLED";
    FD1P3IX SLO__i10 (.D(SLO[8]), .SP(clk_enable_1057), .CD(GND_net), 
            .CK(clk), .Q(SLO[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i10.GSR = "DISABLED";
    FD1P3IX SLO__i14 (.D(SLO[12]), .SP(clk_enable_1057), .CD(GND_net), 
            .CK(clk), .Q(SLO[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i14.GSR = "DISABLED";
    FD1P3IX SLO__i17 (.D(SLO[15]), .SP(clk_enable_1057), .CD(GND_net), 
            .CK(clk), .Q(SLO[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i17.GSR = "DISABLED";
    FD1P3IX SLO__i11 (.D(SLO[9]), .SP(clk_enable_1057), .CD(GND_net), 
            .CK(clk), .Q(SLO[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i11.GSR = "DISABLED";
    FD1P3IX SLO__i15 (.D(SLO[13]), .SP(clk_enable_1057), .CD(GND_net), 
            .CK(clk), .Q(SLO[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i15.GSR = "DISABLED";
    FD1P3IX SLO__i18 (.D(SLO[16]), .SP(clk_enable_1057), .CD(GND_net), 
            .CK(clk), .Q(SLO[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i18.GSR = "DISABLED";
    FD1P3IX SLO__i8 (.D(SLO[6]), .SP(clk_enable_1057), .CD(GND_net), .CK(clk), 
            .Q(SLO[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i8.GSR = "DISABLED";
    FD1P3IX SLO__i12 (.D(SLO[10]), .SP(clk_enable_1057), .CD(GND_net), 
            .CK(clk), .Q(SLO[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i12.GSR = "DISABLED";
    FD1P3IX SLO__i9 (.D(SLO[7]), .SP(clk_enable_1057), .CD(GND_net), .CK(clk), 
            .Q(SLO[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i9.GSR = "DISABLED";
    FD1P3IX SLO__i13 (.D(SLO[11]), .SP(clk_enable_1057), .CD(GND_net), 
            .CK(clk), .Q(SLO[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i13.GSR = "DISABLED";
    FD1P3IX SLO__i16 (.D(SLO[14]), .SP(clk_enable_1057), .CD(GND_net), 
            .CK(clk), .Q(SLO[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i16.GSR = "DISABLED";
    FD1P3IX SLO__i19 (.D(SLO[17]), .SP(clk_enable_1057), .CD(GND_net), 
            .CK(clk), .Q(SLO[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i19.GSR = "DISABLED";
    FD1P3IX SLO__i2 (.D(SLO[0]), .SP(clk_enable_1057), .CD(GND_net), .CK(clk), 
            .Q(SLO[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i2.GSR = "DISABLED";
    FD1P3IX SLO__i5 (.D(SLO[3]), .SP(clk_enable_1057), .CD(GND_net), .CK(clk), 
            .Q(SLO[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i5.GSR = "DISABLED";
    FD1P3IX SLO__i3 (.D(SLO[1]), .SP(clk_enable_1057), .CD(GND_net), .CK(clk), 
            .Q(SLO[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i3.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_711 (.A(mode[0]), .B(mode[1]), .Z(n30111)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_rep_711.init = 16'heeee;
    LUT4 i1_2_lut_rep_647_3_lut (.A(mode[0]), .B(mode[1]), .C(mode[2]), 
         .Z(n30047)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_rep_647_3_lut.init = 16'hefef;
    FD1P3IX SLO__i6 (.D(SLO[4]), .SP(clk_enable_1057), .CD(GND_net), .CK(clk), 
            .Q(SLO[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i6.GSR = "DISABLED";
    FD1P3IX SLO__i4 (.D(SLO[2]), .SP(clk_enable_1057), .CD(GND_net), .CK(clk), 
            .Q(SLO[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i4.GSR = "DISABLED";
    FD1P3IX SLO__i7 (.D(SLO[5]), .SP(clk_enable_1057), .CD(GND_net), .CK(clk), 
            .Q(SLO[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i7.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(mode[0]), .B(mode[1]), .C(Cnt[5]), .D(mode[2]), 
         .Z(n26309)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfeff;
    LUT4 i1_2_lut_rep_687_3_lut (.A(mode[0]), .B(mode[1]), .C(mode[2]), 
         .Z(n30087)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_rep_687_3_lut.init = 16'hfefe;
    LUT4 i2991_2_lut_3_lut_4_lut (.A(mode[0]), .B(mode[1]), .C(pin_io_c_54), 
         .D(mode[2]), .Z(\pin_intrpt[17] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2991_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2948_1_lut_2_lut_3_lut (.A(mode[0]), .B(mode[1]), .C(mode[2]), 
         .Z(n7262)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2948_1_lut_2_lut_3_lut.init = 16'h0101;
    LUT4 i2989_2_lut_3_lut_4_lut (.A(mode[0]), .B(mode[1]), .C(pin_io_c_52), 
         .D(mode[2]), .Z(\pin_intrpt[15] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2989_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2990_2_lut_3_lut_4_lut (.A(mode[0]), .B(mode[1]), .C(pin_io_c_53), 
         .D(mode[2]), .Z(\pin_intrpt[16] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2990_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2430_2_lut_rep_712 (.A(mode[0]), .B(mode[1]), .Z(n30112)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2430_2_lut_rep_712.init = 16'h8888;
    LUT4 i24091_2_lut_3_lut (.A(mode[0]), .B(mode[1]), .C(mode[2]), .Z(ENC_O_N_5841)) /* synthesis lut_function=(!(A (B+(C))+!A (C))) */ ;
    defparam i24091_2_lut_3_lut.init = 16'h0707;
    FD1P3AX NSL_484 (.D(NSL_N_5872), .SP(clk_1MHz_enable_69), .CK(clk_1MHz), 
            .Q(NSL)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam NSL_484.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_715 (.A(Cnt[7]), .B(Cnt[6]), .Z(n30115)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(109[8:17])
    defparam i1_2_lut_rep_715.init = 16'heeee;
    LUT4 i1_3_lut_rep_666_4_lut (.A(Cnt[7]), .B(Cnt[6]), .C(Cnt[0]), .D(n30116), 
         .Z(n30066)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(109[8:17])
    defparam i1_3_lut_rep_666_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_716 (.A(Cnt[2]), .B(Cnt[3]), .Z(n30116)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(109[8:17])
    defparam i1_2_lut_rep_716.init = 16'heeee;
    LUT4 i1_3_lut_4_lut (.A(Cnt[2]), .B(Cnt[3]), .C(Cnt[1]), .D(Cnt[0]), 
         .Z(n18446)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(109[8:17])
    defparam i1_3_lut_4_lut.init = 16'hfeee;
    LUT4 i1_3_lut_rep_732 (.A(Cnt_NSL[9]), .B(Cnt_NSL[8]), .C(Cnt_NSL[7]), 
         .Z(n30132)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_rep_732.init = 16'hfefe;
    LUT4 i1_2_lut_rep_657_4_lut (.A(Cnt_NSL[9]), .B(Cnt_NSL[8]), .C(Cnt_NSL[7]), 
         .D(n30133), .Z(n30057)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_rep_657_4_lut.init = 16'hfe00;
    LUT4 i1_2_lut_rep_733 (.A(Cnt_NSL[11]), .B(Cnt_NSL[10]), .Z(n30133)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i1_2_lut_rep_733.init = 16'h8888;
    LUT4 i23937_2_lut_rep_621_3_lut_4_lut (.A(Cnt_NSL[11]), .B(Cnt_NSL[10]), 
         .C(resetn_c), .D(n30132), .Z(clk_1MHz_enable_34)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i23937_2_lut_rep_621_3_lut_4_lut.init = 16'h8f0f;
    LUT4 i23996_2_lut_rep_749 (.A(MA_Temp), .B(clk_1MHz), .Z(n30149)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i23996_2_lut_rep_749.init = 16'h7777;
    LUT4 i1_2_lut_rep_667_3_lut (.A(MA_Temp), .B(clk_1MHz), .C(prev_MA), 
         .Z(n30067)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i1_2_lut_rep_667_3_lut.init = 16'hf8f8;
    
endmodule
//
// Verilog Description of module \io(UART_ADDRESS_WIDTH=4) 
//

module \io(UART_ADDRESS_WIDTH=4)  (pwm_out_1, clk_100k, clk_100k_enable_1, 
            n2193, clk, clk_enable_695, n30185, \spi_data_r[0] , mode, 
            clk_enable_235, \spi_data_r[1] , \spi_data_r[3] , \spi_data_r[4] , 
            \spi_data_r[7] , \spi_data_r[8] , \spi_data_r[9] , \spi_data_r[10] , 
            \spi_data_r[11] , GND_net, pwm_out_1_N_6306, clk_enable_959, 
            \spi_data_r[2] , \spi_data_r[5] , \spi_data_r[6] , n18, 
            resetn_c) /* synthesis syn_module_defined=1 */ ;
    output pwm_out_1;
    input clk_100k;
    input clk_100k_enable_1;
    input n2193;
    input clk;
    input clk_enable_695;
    input n30185;
    input \spi_data_r[0] ;
    output mode;
    input clk_enable_235;
    input \spi_data_r[1] ;
    input \spi_data_r[3] ;
    input \spi_data_r[4] ;
    input \spi_data_r[7] ;
    input \spi_data_r[8] ;
    input \spi_data_r[9] ;
    input \spi_data_r[10] ;
    input \spi_data_r[11] ;
    input GND_net;
    output pwm_out_1_N_6306;
    input clk_enable_959;
    input \spi_data_r[2] ;
    input \spi_data_r[5] ;
    input \spi_data_r[6] ;
    output n18;
    input resetn_c;
    
    wire clk_100k /* synthesis SET_AS_NETWORK=clk_100k, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(134[6:14])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    
    wire n25107;
    wire [11:0]pwm_freq_cntr;   // c:/s_links/sources/slot_cards/slider_io.v(55[33:46])
    wire [11:0]n53;
    wire [11:0]pwm_duty_1;   // c:/s_links/sources/slot_cards/slider_io.v(51[33:43])
    
    wire n21969;
    wire [12:0]pwm_out_1_N_6307;
    
    wire n21968, n21967, n21966, n21965, n21964, n21896, n21895, 
        n21894, n21893, n21892, n21891, n21785, n21784, n21783, 
        n21782, n21, n22, n20, n14, n28376, n27347, n27345, 
        n27335;
    
    FD1P3AX pwm_out_1_130 (.D(n25107), .SP(clk_100k_enable_1), .CK(clk_100k), 
            .Q(pwm_out_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=454, LSE_RLINE=486 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(114[8] 162[4])
    defparam pwm_out_1_130.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1785__i0 (.D(n53[0]), .CK(clk_100k), .CD(n2193), 
            .Q(pwm_freq_cntr[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785__i0.GSR = "DISABLED";
    FD1P3IX pwm_duty_1_i0 (.D(\spi_data_r[0] ), .SP(clk_enable_695), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=454, LSE_RLINE=486 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(94[8] 111[4])
    defparam pwm_duty_1_i0.GSR = "DISABLED";
    FD1P3IX mode_125 (.D(\spi_data_r[0] ), .SP(clk_enable_235), .CD(n30185), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=454, LSE_RLINE=486 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(78[8] 86[4])
    defparam mode_125.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1785__i11 (.D(n53[11]), .CK(clk_100k), .CD(n2193), 
            .Q(pwm_freq_cntr[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785__i11.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1785__i10 (.D(n53[10]), .CK(clk_100k), .CD(n2193), 
            .Q(pwm_freq_cntr[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785__i10.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1785__i9 (.D(n53[9]), .CK(clk_100k), .CD(n2193), 
            .Q(pwm_freq_cntr[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785__i9.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1785__i8 (.D(n53[8]), .CK(clk_100k), .CD(n2193), 
            .Q(pwm_freq_cntr[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785__i8.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1785__i7 (.D(n53[7]), .CK(clk_100k), .CD(n2193), 
            .Q(pwm_freq_cntr[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785__i7.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1785__i6 (.D(n53[6]), .CK(clk_100k), .CD(n2193), 
            .Q(pwm_freq_cntr[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785__i6.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1785__i5 (.D(n53[5]), .CK(clk_100k), .CD(n2193), 
            .Q(pwm_freq_cntr[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785__i5.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1785__i4 (.D(n53[4]), .CK(clk_100k), .CD(n2193), 
            .Q(pwm_freq_cntr[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785__i4.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1785__i3 (.D(n53[3]), .CK(clk_100k), .CD(n2193), 
            .Q(pwm_freq_cntr[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785__i3.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1785__i2 (.D(n53[2]), .CK(clk_100k), .CD(n2193), 
            .Q(pwm_freq_cntr[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785__i2.GSR = "DISABLED";
    FD1S3IX pwm_freq_cntr_1785__i1 (.D(n53[1]), .CK(clk_100k), .CD(n2193), 
            .Q(pwm_freq_cntr[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785__i1.GSR = "DISABLED";
    FD1P3IX pwm_duty_1_i1 (.D(\spi_data_r[1] ), .SP(clk_enable_695), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=454, LSE_RLINE=486 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(94[8] 111[4])
    defparam pwm_duty_1_i1.GSR = "DISABLED";
    FD1P3IX pwm_duty_1_i3 (.D(\spi_data_r[3] ), .SP(clk_enable_695), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=454, LSE_RLINE=486 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(94[8] 111[4])
    defparam pwm_duty_1_i3.GSR = "DISABLED";
    FD1P3IX pwm_duty_1_i4 (.D(\spi_data_r[4] ), .SP(clk_enable_695), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=454, LSE_RLINE=486 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(94[8] 111[4])
    defparam pwm_duty_1_i4.GSR = "DISABLED";
    FD1P3IX pwm_duty_1_i7 (.D(\spi_data_r[7] ), .SP(clk_enable_695), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=454, LSE_RLINE=486 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(94[8] 111[4])
    defparam pwm_duty_1_i7.GSR = "DISABLED";
    FD1P3IX pwm_duty_1_i8 (.D(\spi_data_r[8] ), .SP(clk_enable_695), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=454, LSE_RLINE=486 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(94[8] 111[4])
    defparam pwm_duty_1_i8.GSR = "DISABLED";
    FD1P3IX pwm_duty_1_i9 (.D(\spi_data_r[9] ), .SP(clk_enable_695), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=454, LSE_RLINE=486 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(94[8] 111[4])
    defparam pwm_duty_1_i9.GSR = "DISABLED";
    FD1P3IX pwm_duty_1_i10 (.D(\spi_data_r[10] ), .SP(clk_enable_695), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=454, LSE_RLINE=486 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(94[8] 111[4])
    defparam pwm_duty_1_i10.GSR = "DISABLED";
    FD1P3IX pwm_duty_1_i11 (.D(\spi_data_r[11] ), .SP(clk_enable_695), .CD(n30185), 
            .CK(clk), .Q(pwm_duty_1[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=454, LSE_RLINE=486 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(94[8] 111[4])
    defparam pwm_duty_1_i11.GSR = "DISABLED";
    CCU2D sub_96_add_2_13 (.A0(pwm_duty_1[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21969), .S0(pwm_out_1_N_6307[11]), .S1(pwm_out_1_N_6307[12]));   // c:/s_links/sources/slot_cards/slider_io.v(141[25:39])
    defparam sub_96_add_2_13.INIT0 = 16'h5555;
    defparam sub_96_add_2_13.INIT1 = 16'hffff;
    defparam sub_96_add_2_13.INJECT1_0 = "NO";
    defparam sub_96_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_96_add_2_11 (.A0(pwm_duty_1[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_1[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21968), .COUT(n21969), .S0(pwm_out_1_N_6307[9]), 
          .S1(pwm_out_1_N_6307[10]));   // c:/s_links/sources/slot_cards/slider_io.v(141[25:39])
    defparam sub_96_add_2_11.INIT0 = 16'h5555;
    defparam sub_96_add_2_11.INIT1 = 16'h5555;
    defparam sub_96_add_2_11.INJECT1_0 = "NO";
    defparam sub_96_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_96_add_2_9 (.A0(pwm_duty_1[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_1[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21967), .COUT(n21968), .S0(pwm_out_1_N_6307[7]), 
          .S1(pwm_out_1_N_6307[8]));   // c:/s_links/sources/slot_cards/slider_io.v(141[25:39])
    defparam sub_96_add_2_9.INIT0 = 16'h5555;
    defparam sub_96_add_2_9.INIT1 = 16'h5555;
    defparam sub_96_add_2_9.INJECT1_0 = "NO";
    defparam sub_96_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_96_add_2_7 (.A0(pwm_duty_1[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_1[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21966), .COUT(n21967), .S0(pwm_out_1_N_6307[5]), 
          .S1(pwm_out_1_N_6307[6]));   // c:/s_links/sources/slot_cards/slider_io.v(141[25:39])
    defparam sub_96_add_2_7.INIT0 = 16'h5555;
    defparam sub_96_add_2_7.INIT1 = 16'h5555;
    defparam sub_96_add_2_7.INJECT1_0 = "NO";
    defparam sub_96_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_96_add_2_5 (.A0(pwm_duty_1[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_1[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21965), .COUT(n21966), .S0(pwm_out_1_N_6307[3]), 
          .S1(pwm_out_1_N_6307[4]));   // c:/s_links/sources/slot_cards/slider_io.v(141[25:39])
    defparam sub_96_add_2_5.INIT0 = 16'h5555;
    defparam sub_96_add_2_5.INIT1 = 16'h5555;
    defparam sub_96_add_2_5.INJECT1_0 = "NO";
    defparam sub_96_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_96_add_2_3 (.A0(pwm_duty_1[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty_1[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21964), .COUT(n21965), .S0(pwm_out_1_N_6307[1]), 
          .S1(pwm_out_1_N_6307[2]));   // c:/s_links/sources/slot_cards/slider_io.v(141[25:39])
    defparam sub_96_add_2_3.INIT0 = 16'h5555;
    defparam sub_96_add_2_3.INIT1 = 16'h5555;
    defparam sub_96_add_2_3.INJECT1_0 = "NO";
    defparam sub_96_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_96_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_duty_1[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n21964), .S1(pwm_out_1_N_6307[0]));   // c:/s_links/sources/slot_cards/slider_io.v(141[25:39])
    defparam sub_96_add_2_1.INIT0 = 16'hF000;
    defparam sub_96_add_2_1.INIT1 = 16'h5555;
    defparam sub_96_add_2_1.INJECT1_0 = "NO";
    defparam sub_96_add_2_1.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1785_add_4_13 (.A0(pwm_freq_cntr[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21896), .S0(n53[11]));   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785_add_4_13.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1785_add_4_13.INIT1 = 16'h0000;
    defparam pwm_freq_cntr_1785_add_4_13.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1785_add_4_13.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1785_add_4_11 (.A0(pwm_freq_cntr[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n21895), .COUT(n21896), .S0(n53[9]), 
          .S1(n53[10]));   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785_add_4_11.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1785_add_4_11.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1785_add_4_11.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1785_add_4_11.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1785_add_4_9 (.A0(pwm_freq_cntr[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n21894), .COUT(n21895), .S0(n53[7]), 
          .S1(n53[8]));   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785_add_4_9.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1785_add_4_9.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1785_add_4_9.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1785_add_4_9.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1785_add_4_7 (.A0(pwm_freq_cntr[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n21893), .COUT(n21894), .S0(n53[5]), 
          .S1(n53[6]));   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785_add_4_7.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1785_add_4_7.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1785_add_4_7.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1785_add_4_7.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1785_add_4_5 (.A0(pwm_freq_cntr[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n21892), .COUT(n21893), .S0(n53[3]), 
          .S1(n53[4]));   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785_add_4_5.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1785_add_4_5.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1785_add_4_5.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1785_add_4_5.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1785_add_4_3 (.A0(pwm_freq_cntr[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n21891), .COUT(n21892), .S0(n53[1]), 
          .S1(n53[2]));   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785_add_4_3.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_1785_add_4_3.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_1785_add_4_3.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1785_add_4_3.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_1785_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_freq_cntr[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n21891), .S1(n53[0]));   // c:/s_links/sources/slot_cards/slider_io.v(159[22:42])
    defparam pwm_freq_cntr_1785_add_4_1.INIT0 = 16'hF000;
    defparam pwm_freq_cntr_1785_add_4_1.INIT1 = 16'h0555;
    defparam pwm_freq_cntr_1785_add_4_1.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_1785_add_4_1.INJECT1_1 = "NO";
    CCU2D equal_180_13 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21785), 
          .S0(pwm_out_1_N_6306));
    defparam equal_180_13.INIT0 = 16'hFFFF;
    defparam equal_180_13.INIT1 = 16'h0000;
    defparam equal_180_13.INJECT1_0 = "NO";
    defparam equal_180_13.INJECT1_1 = "NO";
    CCU2D equal_180_13_17467 (.A0(pwm_out_1_N_6307[3]), .B0(pwm_freq_cntr[3]), 
          .C0(pwm_out_1_N_6307[2]), .D0(pwm_freq_cntr[2]), .A1(pwm_out_1_N_6307[1]), 
          .B1(pwm_freq_cntr[1]), .C1(pwm_out_1_N_6307[0]), .D1(pwm_freq_cntr[0]), 
          .CIN(n21784), .COUT(n21785));
    defparam equal_180_13_17467.INIT0 = 16'h9009;
    defparam equal_180_13_17467.INIT1 = 16'h9009;
    defparam equal_180_13_17467.INJECT1_0 = "YES";
    defparam equal_180_13_17467.INJECT1_1 = "YES";
    CCU2D equal_180_11 (.A0(pwm_out_1_N_6307[7]), .B0(pwm_freq_cntr[7]), 
          .C0(pwm_out_1_N_6307[6]), .D0(pwm_freq_cntr[6]), .A1(pwm_out_1_N_6307[5]), 
          .B1(pwm_freq_cntr[5]), .C1(pwm_out_1_N_6307[4]), .D1(pwm_freq_cntr[4]), 
          .CIN(n21783), .COUT(n21784));
    defparam equal_180_11.INIT0 = 16'h9009;
    defparam equal_180_11.INIT1 = 16'h9009;
    defparam equal_180_11.INJECT1_0 = "YES";
    defparam equal_180_11.INJECT1_1 = "YES";
    CCU2D equal_180_9 (.A0(pwm_out_1_N_6307[11]), .B0(pwm_freq_cntr[11]), 
          .C0(pwm_out_1_N_6307[10]), .D0(pwm_freq_cntr[10]), .A1(pwm_out_1_N_6307[9]), 
          .B1(pwm_freq_cntr[9]), .C1(pwm_out_1_N_6307[8]), .D1(pwm_freq_cntr[8]), 
          .CIN(n21782), .COUT(n21783));
    defparam equal_180_9.INIT0 = 16'h9009;
    defparam equal_180_9.INIT1 = 16'h9009;
    defparam equal_180_9.INJECT1_0 = "YES";
    defparam equal_180_9.INJECT1_1 = "YES";
    CCU2D equal_180_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_out_1_N_6307[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n21782));   // c:/s_links/sources/slot_cards/slider_io.v(141[8:39])
    defparam equal_180_0.INIT0 = 16'hF000;
    defparam equal_180_0.INIT1 = 16'h5555;
    defparam equal_180_0.INJECT1_0 = "NO";
    defparam equal_180_0.INJECT1_1 = "YES";
    FD1P3JX pwm_duty_1_i2 (.D(\spi_data_r[2] ), .SP(clk_enable_959), .PD(n30185), 
            .CK(clk), .Q(pwm_duty_1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=454, LSE_RLINE=486 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(94[8] 111[4])
    defparam pwm_duty_1_i2.GSR = "DISABLED";
    FD1P3JX pwm_duty_1_i5 (.D(\spi_data_r[5] ), .SP(clk_enable_959), .PD(n30185), 
            .CK(clk), .Q(pwm_duty_1[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=454, LSE_RLINE=486 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(94[8] 111[4])
    defparam pwm_duty_1_i5.GSR = "DISABLED";
    FD1P3JX pwm_duty_1_i6 (.D(\spi_data_r[6] ), .SP(clk_enable_959), .PD(n30185), 
            .CK(clk), .Q(pwm_duty_1[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=454, LSE_RLINE=486 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(94[8] 111[4])
    defparam pwm_duty_1_i6.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(n21), .B(n18), .C(resetn_c), .D(n22), .Z(n25107)) /* synthesis lut_function=(A (B (C))+!A (B (C (D)))) */ ;   // c:/s_links/sources/mcm_top.v(17[27:33])
    defparam i1_4_lut.init = 16'hc080;
    LUT4 i9_4_lut (.A(pwm_duty_1[7]), .B(pwm_duty_1[9]), .C(pwm_duty_1[6]), 
         .D(pwm_duty_1[4]), .Z(n21)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/slider_io.v(51[33:43])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i10_4_lut (.A(pwm_duty_1[1]), .B(n20), .C(n14), .D(pwm_duty_1[2]), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/slider_io.v(51[33:43])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i8_4_lut (.A(pwm_duty_1[10]), .B(pwm_duty_1[11]), .C(pwm_duty_1[0]), 
         .D(pwm_duty_1[5]), .Z(n20)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/slider_io.v(51[33:43])
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(pwm_duty_1[3]), .B(pwm_duty_1[8]), .Z(n14)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/slider_io.v(51[33:43])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_844 (.A(n28376), .B(pwm_freq_cntr[4]), .C(n27347), 
         .D(n27345), .Z(n18)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_844.init = 16'h1000;
    LUT4 i23674_2_lut (.A(pwm_freq_cntr[5]), .B(pwm_freq_cntr[11]), .Z(n28376)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23674_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_845 (.A(pwm_freq_cntr[1]), .B(n27335), .C(pwm_freq_cntr[2]), 
         .D(pwm_freq_cntr[0]), .Z(n27347)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/s_links/sources/mcm_top.v(17[27:33])
    defparam i1_4_lut_adj_845.init = 16'h8000;
    LUT4 i1_4_lut_adj_846 (.A(pwm_freq_cntr[6]), .B(pwm_freq_cntr[8]), .C(pwm_freq_cntr[9]), 
         .D(pwm_freq_cntr[10]), .Z(n27345)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/s_links/sources/mcm_top.v(17[27:33])
    defparam i1_4_lut_adj_846.init = 16'h8000;
    LUT4 i1_2_lut (.A(pwm_freq_cntr[3]), .B(pwm_freq_cntr[7]), .Z(n27335)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/mcm_top.v(17[27:33])
    defparam i1_2_lut.init = 16'h8888;
    
endmodule
//
// Verilog Description of module \stepper(UART_ADDRESS_WIDTH=4) 
//

module \stepper(UART_ADDRESS_WIDTH=4)  (GND_net, clk, \spi_addr_r[0] , 
            n30070, n23526, n30035, n29990, clk_1MHz, n30185, resetn_c, 
            n30129, spi_data_out_r_39__N_3825, pin_io_out_8, spi_data_out_r_39__N_3865, 
            mode_adj_654, clk_enable_761, \spi_data_r[0] , n30175, n30058, 
            digital_output_r, n28547, n47, \spi_addr_r[1] , n26957, 
            n23537, n20647, n23978, \spi_cmd_r[2] , \spi_cmd_r[8] , 
            \spi_cmd_r[10] , \spi_cmd_r[6] , \spi_cmd_r[7] , \spi_cmd_r[12] , 
            \spi_cmd_r[15] , n30134, n30125, mode, n23609, n30138, 
            n23916, n25979, clk_enable_222, n26633, n30028, n26779, 
            n30198, n32, \spi_data_r[1] , \spi_data_r[2] , NSL, EM_STOP, 
            n25721, n25547, n24169, n18440, n28402, n28524, n30045, 
            n29999, n28486, \spi_addr_r[4] , \spi_addr_r[2] , n27013, 
            \spi_cmd_r[0] , spi_data_valid_r, \spi_addr_r[3] , n30052, 
            n30007, clk_enable_242, n29994, n30199, n25739, n25699, 
            n25941, n25943, n25801, \spi_cmd_r[3] , n30044, clk_enable_256, 
            \spi_cmd_r[1] , \spi_cmd_r[4] , \spi_cmd_r[5] , reset_r, 
            reset_r_N_4129, n30043, mode_adj_653, n30018, pin_io_out_4, 
            \pin_intrpt[2] , \quad_homing[0] , n25869, n30151) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk;
    input \spi_addr_r[0] ;
    input n30070;
    input n23526;
    input n30035;
    output n29990;
    input clk_1MHz;
    input n30185;
    input resetn_c;
    output n30129;
    output [39:0]spi_data_out_r_39__N_3825;
    input pin_io_out_8;
    output spi_data_out_r_39__N_3865;
    output [2:0]mode_adj_654;
    input clk_enable_761;
    input \spi_data_r[0] ;
    output n30175;
    output n30058;
    output digital_output_r;
    input n28547;
    input n47;
    input \spi_addr_r[1] ;
    output n26957;
    input n23537;
    output n20647;
    input n23978;
    input \spi_cmd_r[2] ;
    input \spi_cmd_r[8] ;
    input \spi_cmd_r[10] ;
    input \spi_cmd_r[6] ;
    input \spi_cmd_r[7] ;
    input \spi_cmd_r[12] ;
    input \spi_cmd_r[15] ;
    output n30134;
    input n30125;
    input mode;
    output n23609;
    input n30138;
    input n23916;
    input n25979;
    output clk_enable_222;
    input n26633;
    output n30028;
    input n26779;
    input n30198;
    input n32;
    input \spi_data_r[1] ;
    input \spi_data_r[2] ;
    output NSL;
    input EM_STOP;
    input n25721;
    input n25547;
    output n24169;
    output n18440;
    input n28402;
    input n28524;
    output n30045;
    output n29999;
    input n28486;
    input \spi_addr_r[4] ;
    input \spi_addr_r[2] ;
    output n27013;
    input \spi_cmd_r[0] ;
    input spi_data_valid_r;
    input \spi_addr_r[3] ;
    output n30052;
    output n30007;
    output clk_enable_242;
    output n29994;
    output n30199;
    input n25739;
    output n25699;
    input n25941;
    output n25943;
    output n25801;
    input \spi_cmd_r[3] ;
    input n30044;
    output clk_enable_256;
    input \spi_cmd_r[1] ;
    input \spi_cmd_r[4] ;
    input \spi_cmd_r[5] ;
    output reset_r;
    input reset_r_N_4129;
    output n30043;
    input mode_adj_653;
    output n30018;
    input pin_io_out_4;
    output \pin_intrpt[2] ;
    input \quad_homing[0] ;
    output n25869;
    output n30151;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire clk_1MHz /* synthesis SET_AS_NETWORK=clk_1MHz, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(136[6:14])
    wire \pin_intrpt[2]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[2] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    
    wire n21915;
    wire [7:0]Cnt;   // c:/s_links/sources/slot_cards/stepper.v(62[11:14])
    wire [31:0]n153;
    
    wire n21916;
    wire [51:0]SLO;   // c:/s_links/sources/slot_cards/stepper.v(63[12:15])
    
    wire clk_enable_1132, n12235;
    wire [51:0]SLO_buf;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire SLO_buf_51__N_4015, MA_Temp, clk_1MHz_enable_7, MA_Temp_N_4144;
    wire [11:0]n93;
    wire [11:0]n53;
    
    wire prev_MA_Temp, n21914, prev_MA;
    wire [39:0]spi_data_out_r_39__N_4076;
    
    wire spi_data_out_r_39__N_4162, clk_1MHz_enable_56;
    wire [7:0]n199;
    
    wire n30130, n24814, n18584, n30077, n18404, n18522, clk_enable_212, 
        n30109, n30172, n25487, n28414, n28504, n28420, n25471, 
        n26363, n30063;
    wire [11:0]Cnt_NSL;   // c:/s_links/sources/slot_cards/stepper.v(61[12:19])
    
    wire n28585, n28586, n21906, n21905, n30078, n30005, NSL_N_4157, 
        clk_enable_1104, n21904, n21903, n4, n28326, n30056, n21902, 
        n30131, n30177, n30176, clk_1MHz_enable_65, n21901, n30190, 
        n25793, n21917;
    
    CCU2D add_564_5 (.A0(Cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21915), 
          .COUT(n21916), .S0(n153[3]), .S1(n153[4]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_5.INIT0 = 16'h5aaa;
    defparam add_564_5.INIT1 = 16'h5aaa;
    defparam add_564_5.INJECT1_0 = "NO";
    defparam add_564_5.INJECT1_1 = "NO";
    FD1P3IX SLO__i42 (.D(SLO[40]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i42.GSR = "DISABLED";
    FD1P3AX SLO_buf__i1 (.D(SLO[0]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i1.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_590_3_lut_4_lut (.A(\spi_addr_r[0] ), .B(n30070), 
         .C(n23526), .D(n30035), .Z(n29990)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_rep_590_3_lut_4_lut.init = 16'h2000;
    FD1P3IX MA_Temp_483 (.D(MA_Temp_N_4144), .SP(clk_1MHz_enable_7), .CD(n30185), 
            .CK(clk_1MHz), .Q(MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam MA_Temp_483.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1778__i0 (.D(n53[0]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778__i0.GSR = "DISABLED";
    FD1P3IX SLO__i43 (.D(SLO[41]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i43.GSR = "DISABLED";
    FD1S3AX prev_MA_Temp_487 (.D(MA_Temp), .CK(clk), .Q(prev_MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam prev_MA_Temp_487.GSR = "DISABLED";
    CCU2D add_564_3 (.A0(Cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21914), 
          .COUT(n21915), .S0(n153[1]), .S1(n153[2]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_3.INIT0 = 16'h5aaa;
    defparam add_564_3.INIT1 = 16'h5aaa;
    defparam add_564_3.INJECT1_0 = "NO";
    defparam add_564_3.INJECT1_1 = "NO";
    FD1S3AX prev_MA_489 (.D(n30129), .CK(clk), .Q(prev_MA)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam prev_MA_489.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i0 (.D(spi_data_out_r_39__N_4076[0]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i0.GSR = "DISABLED";
    FD1P3IX SLO__i1 (.D(pin_io_out_8), .SP(clk_enable_1132), .CD(GND_net), 
            .CK(clk), .Q(SLO[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i1.GSR = "DISABLED";
    CCU2D add_564_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n21914), 
          .S1(n153[0]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_1.INIT0 = 16'hF000;
    defparam add_564_1.INIT1 = 16'h5555;
    defparam add_564_1.INJECT1_0 = "NO";
    defparam add_564_1.INJECT1_1 = "NO";
    FD1P3IX SLO__i2 (.D(SLO[0]), .SP(clk_enable_1132), .CD(GND_net), .CK(clk), 
            .Q(SLO[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i2.GSR = "DISABLED";
    FD1P3IX SLO__i3 (.D(SLO[1]), .SP(clk_enable_1132), .CD(GND_net), .CK(clk), 
            .Q(SLO[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i3.GSR = "DISABLED";
    FD1S3IX i168_494 (.D(spi_data_out_r_39__N_4162), .CK(clk), .CD(n30185), 
            .Q(spi_data_out_r_39__N_3865)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam i168_494.GSR = "DISABLED";
    FD1P3IX SLO__i4 (.D(SLO[2]), .SP(clk_enable_1132), .CD(GND_net), .CK(clk), 
            .Q(SLO[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i4.GSR = "DISABLED";
    FD1P3IX SLO__i5 (.D(SLO[3]), .SP(clk_enable_1132), .CD(GND_net), .CK(clk), 
            .Q(SLO[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i5.GSR = "DISABLED";
    FD1P3IX SLO__i6 (.D(SLO[4]), .SP(clk_enable_1132), .CD(GND_net), .CK(clk), 
            .Q(SLO[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i6.GSR = "DISABLED";
    FD1P3IX SLO__i7 (.D(SLO[5]), .SP(clk_enable_1132), .CD(GND_net), .CK(clk), 
            .Q(SLO[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i7.GSR = "DISABLED";
    FD1P3IX Cnt__i0 (.D(n199[0]), .SP(clk_1MHz_enable_56), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i0.GSR = "DISABLED";
    FD1P3IX SLO__i44 (.D(SLO[42]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i44.GSR = "DISABLED";
    FD1P3IX mode__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_761), .CD(n30185), 
            .CK(clk), .Q(mode_adj_654[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i0.GSR = "DISABLED";
    FD1P3IX SLO__i8 (.D(SLO[6]), .SP(clk_enable_1132), .CD(GND_net), .CK(clk), 
            .Q(SLO[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i8.GSR = "DISABLED";
    FD1P3IX SLO__i45 (.D(SLO[43]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i45.GSR = "DISABLED";
    FD1P3IX SLO__i46 (.D(SLO[44]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i46.GSR = "DISABLED";
    FD1P3IX SLO__i9 (.D(SLO[7]), .SP(clk_enable_1132), .CD(GND_net), .CK(clk), 
            .Q(SLO[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i9.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(n30130), .B(n24814), .C(n30175), .D(mode_adj_654[2]), 
         .Z(n18584)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(107[27:54])
    defparam i1_4_lut.init = 16'hffef;
    LUT4 i1_3_lut (.A(Cnt[5]), .B(n30077), .C(Cnt[4]), .Z(n24814)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_adj_831 (.A(n30130), .B(n18404), .C(Cnt[5]), .D(n30058), 
         .Z(n18522)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam i1_4_lut_adj_831.init = 16'hfffe;
    FD1P3IX digital_output_r_492 (.D(n28547), .SP(clk_enable_212), .CD(n30185), 
            .CK(clk), .Q(digital_output_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam digital_output_r_492.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i39 (.D(SLO_buf[13]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i39.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i38 (.D(SLO_buf[12]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i38.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i37 (.D(SLO_buf[11]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i37.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i36 (.D(SLO_buf[10]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i36.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i35 (.D(spi_data_out_r_39__N_4076[35]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i35.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i34 (.D(spi_data_out_r_39__N_4076[34]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i34.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i33 (.D(spi_data_out_r_39__N_4076[33]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i33.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(spi_data_out_r_39__N_4076[32]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i31 (.D(SLO_buf[45]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i30 (.D(SLO_buf[44]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i29 (.D(SLO_buf[43]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i28 (.D(SLO_buf[42]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i27 (.D(SLO_buf[41]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i26 (.D(SLO_buf[40]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i25 (.D(SLO_buf[39]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i24 (.D(SLO_buf[38]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i23 (.D(SLO_buf[37]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i22 (.D(SLO_buf[36]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i21 (.D(SLO_buf[35]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i20 (.D(SLO_buf[34]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i19 (.D(SLO_buf[33]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i18 (.D(SLO_buf[32]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i17 (.D(SLO_buf[31]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i16 (.D(SLO_buf[30]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_3825[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(spi_data_out_r_39__N_4076[15]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(spi_data_out_r_39__N_4076[14]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(spi_data_out_r_39__N_4076[13]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(spi_data_out_r_39__N_4076[12]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(spi_data_out_r_39__N_4076[11]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(spi_data_out_r_39__N_4076[10]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(spi_data_out_r_39__N_4076[9]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(spi_data_out_r_39__N_4076[8]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(spi_data_out_r_39__N_4076[7]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(spi_data_out_r_39__N_4076[6]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(spi_data_out_r_39__N_4076[5]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(spi_data_out_r_39__N_4076[4]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(spi_data_out_r_39__N_4076[3]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(spi_data_out_r_39__N_4076[2]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(spi_data_out_r_39__N_4076[1]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3825[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut (.A(n30109), .B(\spi_addr_r[1] ), .C(n30172), 
         .D(n30070), .Z(n26957)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0010;
    FD1P3IX SLO__i10 (.D(SLO[8]), .SP(clk_enable_1132), .CD(GND_net), 
            .CK(clk), .Q(SLO[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i10.GSR = "DISABLED";
    FD1P3IX SLO__i11 (.D(SLO[9]), .SP(clk_enable_1132), .CD(GND_net), 
            .CK(clk), .Q(SLO[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i11.GSR = "DISABLED";
    FD1P3IX SLO__i12 (.D(SLO[10]), .SP(clk_enable_1132), .CD(GND_net), 
            .CK(clk), .Q(SLO[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i12.GSR = "DISABLED";
    FD1P3IX SLO__i13 (.D(SLO[11]), .SP(clk_enable_1132), .CD(GND_net), 
            .CK(clk), .Q(SLO[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i13.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_832 (.A(n23537), .B(n30070), .C(n25487), .D(n28414), 
         .Z(n20647)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_4_lut_adj_832.init = 16'h0020;
    LUT4 i1_4_lut_adj_833 (.A(n28504), .B(n23978), .C(n28420), .D(n25471), 
         .Z(n25487)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_833.init = 16'h0100;
    LUT4 i23712_2_lut (.A(\spi_cmd_r[2] ), .B(\spi_addr_r[1] ), .Z(n28414)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23712_2_lut.init = 16'heeee;
    LUT4 i23802_4_lut (.A(\spi_cmd_r[8] ), .B(\spi_cmd_r[10] ), .C(\spi_cmd_r[6] ), 
         .D(\spi_cmd_r[7] ), .Z(n28504)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23802_4_lut.init = 16'hfffe;
    LUT4 i23718_2_lut (.A(\spi_cmd_r[12] ), .B(\spi_cmd_r[15] ), .Z(n28420)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23718_2_lut.init = 16'heeee;
    LUT4 i24199_4_lut_4_lut (.A(mode_adj_654[2]), .B(n30134), .C(n26363), 
         .D(n30063), .Z(clk_enable_1132)) /* synthesis lut_function=(!(A (B+(D))+!A ((D)+!C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i24199_4_lut_4_lut.init = 16'h0072;
    LUT4 i24035_2_lut_3_lut_4_lut (.A(mode_adj_654[2]), .B(n30134), .C(n30125), 
         .D(mode), .Z(n23609)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i24035_2_lut_3_lut_4_lut.init = 16'h00d0;
    FD1P3AX Cnt_NSL_1778__i11 (.D(n53[11]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778__i11.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1778__i10 (.D(n53[10]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778__i10.GSR = "DISABLED";
    FD1P3IX SLO__i14 (.D(SLO[12]), .SP(clk_enable_1132), .CD(GND_net), 
            .CK(clk), .Q(SLO[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i14.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1778__i9 (.D(n53[9]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778__i9.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1778__i8 (.D(n53[8]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778__i8.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1778__i7 (.D(n53[7]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778__i7.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1778__i6 (.D(n53[6]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778__i6.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1778__i5 (.D(n53[5]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778__i5.GSR = "DISABLED";
    FD1P3IX SLO__i15 (.D(SLO[13]), .SP(clk_enable_1132), .CD(GND_net), 
            .CK(clk), .Q(SLO[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i15.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1778__i4 (.D(n53[4]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778__i4.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1778__i3 (.D(n53[3]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778__i3.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1778__i2 (.D(n53[2]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778__i2.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1778__i1 (.D(n53[1]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778__i1.GSR = "DISABLED";
    FD1P3IX SLO__i16 (.D(SLO[14]), .SP(clk_enable_1132), .CD(GND_net), 
            .CK(clk), .Q(SLO[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i16.GSR = "DISABLED";
    LUT4 i24011_3_lut_4_lut (.A(\spi_cmd_r[2] ), .B(n30138), .C(n23916), 
         .D(n25979), .Z(clk_enable_222)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i24011_3_lut_4_lut.init = 16'hbfff;
    FD1P3IX SLO__i17 (.D(SLO[15]), .SP(clk_enable_1132), .CD(GND_net), 
            .CK(clk), .Q(SLO[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i17.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_628_4_lut (.A(\spi_cmd_r[2] ), .B(n30138), .C(n23916), 
         .D(n26633), .Z(n30028)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_3_lut_rep_628_4_lut.init = 16'h4000;
    FD1P3IX SLO__i18 (.D(SLO[16]), .SP(clk_enable_1132), .CD(GND_net), 
            .CK(clk), .Q(SLO[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i18.GSR = "DISABLED";
    FD1P3IX SLO__i19 (.D(SLO[17]), .SP(clk_enable_1132), .CD(GND_net), 
            .CK(clk), .Q(SLO[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i19.GSR = "DISABLED";
    FD1P3IX SLO__i20 (.D(SLO[18]), .SP(clk_enable_1132), .CD(GND_net), 
            .CK(clk), .Q(SLO[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i20.GSR = "DISABLED";
    FD1P3IX SLO__i21 (.D(SLO[19]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i21.GSR = "DISABLED";
    FD1P3IX SLO__i22 (.D(SLO[20]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i22.GSR = "DISABLED";
    LUT4 i24132_2_lut_3_lut_4_lut (.A(prev_MA), .B(n30129), .C(n30134), 
         .D(mode_adj_654[2]), .Z(n12235)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i24132_2_lut_3_lut_4_lut.init = 16'h0400;
    FD1P3IX SLO__i23 (.D(SLO[21]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i23.GSR = "DISABLED";
    FD1P3IX SLO__i24 (.D(SLO[22]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i24.GSR = "DISABLED";
    LUT4 mux_158_i1_3_lut (.A(SLO_buf[14]), .B(SLO_buf[4]), .C(n47), .Z(spi_data_out_r_39__N_4076[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i1_3_lut.init = 16'hcaca;
    FD1P3AX SLO_buf__i46 (.D(SLO[45]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i46.GSR = "DISABLED";
    FD1P3AX SLO_buf__i45 (.D(SLO[44]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i45.GSR = "DISABLED";
    FD1P3AX SLO_buf__i44 (.D(SLO[43]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i44.GSR = "DISABLED";
    FD1P3AX SLO_buf__i43 (.D(SLO[42]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i43.GSR = "DISABLED";
    FD1P3AX SLO_buf__i42 (.D(SLO[41]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i42.GSR = "DISABLED";
    FD1P3AX SLO_buf__i41 (.D(SLO[40]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i41.GSR = "DISABLED";
    FD1P3AX SLO_buf__i40 (.D(SLO[39]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i40.GSR = "DISABLED";
    FD1P3AX SLO_buf__i39 (.D(SLO[38]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i39.GSR = "DISABLED";
    FD1P3AX SLO_buf__i38 (.D(SLO[37]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i38.GSR = "DISABLED";
    FD1P3AX SLO_buf__i37 (.D(SLO[36]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i37.GSR = "DISABLED";
    FD1P3AX SLO_buf__i36 (.D(SLO[35]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i36.GSR = "DISABLED";
    FD1P3AX SLO_buf__i35 (.D(SLO[34]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i35.GSR = "DISABLED";
    FD1P3AX SLO_buf__i34 (.D(SLO[33]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i34.GSR = "DISABLED";
    FD1P3AX SLO_buf__i33 (.D(SLO[32]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i33.GSR = "DISABLED";
    FD1P3AX SLO_buf__i32 (.D(SLO[31]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i32.GSR = "DISABLED";
    FD1P3AX SLO_buf__i31 (.D(SLO[30]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i31.GSR = "DISABLED";
    FD1P3AX SLO_buf__i30 (.D(SLO[29]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i30.GSR = "DISABLED";
    FD1P3AX SLO_buf__i29 (.D(SLO[28]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i29.GSR = "DISABLED";
    FD1P3AX SLO_buf__i28 (.D(SLO[27]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i28.GSR = "DISABLED";
    FD1P3AX SLO_buf__i27 (.D(SLO[26]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i27.GSR = "DISABLED";
    FD1P3AX SLO_buf__i26 (.D(SLO[25]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i26.GSR = "DISABLED";
    FD1P3AX SLO_buf__i25 (.D(SLO[24]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i25.GSR = "DISABLED";
    FD1P3AX SLO_buf__i24 (.D(SLO[23]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i24.GSR = "DISABLED";
    FD1P3AX SLO_buf__i23 (.D(SLO[22]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i23.GSR = "DISABLED";
    FD1P3AX SLO_buf__i22 (.D(SLO[21]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i22.GSR = "DISABLED";
    FD1P3AX SLO_buf__i21 (.D(SLO[20]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i21.GSR = "DISABLED";
    FD1P3AX SLO_buf__i20 (.D(SLO[19]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i20.GSR = "DISABLED";
    FD1P3AX SLO_buf__i19 (.D(SLO[18]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i19.GSR = "DISABLED";
    FD1P3AX SLO_buf__i18 (.D(SLO[17]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i18.GSR = "DISABLED";
    FD1P3AX SLO_buf__i17 (.D(SLO[16]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i17.GSR = "DISABLED";
    FD1P3AX SLO_buf__i16 (.D(SLO[15]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i16.GSR = "DISABLED";
    FD1P3AX SLO_buf__i15 (.D(SLO[14]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i15.GSR = "DISABLED";
    FD1P3AX SLO_buf__i14 (.D(SLO[13]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i14.GSR = "DISABLED";
    FD1P3AX SLO_buf__i13 (.D(SLO[12]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i13.GSR = "DISABLED";
    FD1P3AX SLO_buf__i12 (.D(SLO[11]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i12.GSR = "DISABLED";
    FD1P3AX SLO_buf__i11 (.D(SLO[10]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i11.GSR = "DISABLED";
    FD1P3AX SLO_buf__i10 (.D(SLO[9]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i10.GSR = "DISABLED";
    FD1P3AX SLO_buf__i9 (.D(SLO[8]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i9.GSR = "DISABLED";
    FD1P3AX SLO_buf__i8 (.D(SLO[7]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i8.GSR = "DISABLED";
    FD1P3AX SLO_buf__i7 (.D(SLO[6]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i7.GSR = "DISABLED";
    FD1P3AX SLO_buf__i6 (.D(SLO[5]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i6.GSR = "DISABLED";
    FD1P3AX SLO_buf__i5 (.D(SLO[4]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i5.GSR = "DISABLED";
    FD1P3AX SLO_buf__i4 (.D(SLO[3]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i4.GSR = "DISABLED";
    FD1P3AX SLO_buf__i3 (.D(SLO[2]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i3.GSR = "DISABLED";
    FD1P3AX SLO_buf__i2 (.D(SLO[1]), .SP(SLO_buf_51__N_4015), .CK(clk), 
            .Q(SLO_buf[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i2.GSR = "DISABLED";
    PFUMX MA_Temp_I_109 (.BLUT(n28585), .ALUT(n28586), .C0(n18522), .Z(MA_Temp_N_4144)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;
    LUT4 SLO_buf_51__I_94_2_lut (.A(prev_MA_Temp), .B(MA_Temp), .Z(SLO_buf_51__N_4015)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[5:38])
    defparam SLO_buf_51__I_94_2_lut.init = 16'h2222;
    FD1P3IX SLO__i25 (.D(SLO[23]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i25.GSR = "DISABLED";
    FD1P3IX SLO__i26 (.D(SLO[24]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i26.GSR = "DISABLED";
    FD1P3IX SLO__i27 (.D(SLO[25]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i27.GSR = "DISABLED";
    FD1P3IX SLO__i28 (.D(SLO[26]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i28.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_834 (.A(n47), .B(n26779), .C(n30198), .D(n32), 
         .Z(spi_data_out_r_39__N_4162)) /* synthesis lut_function=(!(A ((C+(D))+!B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(171[15:42])
    defparam i1_4_lut_adj_834.init = 16'h555d;
    FD1P3IX Cnt__i1 (.D(n199[1]), .SP(clk_1MHz_enable_56), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i1.GSR = "DISABLED";
    FD1P3IX Cnt__i2 (.D(n199[2]), .SP(clk_1MHz_enable_56), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i3 (.D(n199[3]), .SP(clk_1MHz_enable_56), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i3.GSR = "DISABLED";
    FD1P3IX Cnt__i4 (.D(n199[4]), .SP(clk_1MHz_enable_56), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i4.GSR = "DISABLED";
    FD1P3IX Cnt__i5 (.D(n199[5]), .SP(clk_1MHz_enable_56), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i5.GSR = "DISABLED";
    FD1P3IX Cnt__i6 (.D(n199[6]), .SP(clk_1MHz_enable_56), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i6.GSR = "DISABLED";
    FD1P3IX Cnt__i7 (.D(n199[7]), .SP(clk_1MHz_enable_56), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i7.GSR = "DISABLED";
    FD1P3IX mode__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_761), .CD(n30185), 
            .CK(clk), .Q(mode_adj_654[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i1.GSR = "DISABLED";
    FD1P3IX mode__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_761), .CD(n30185), 
            .CK(clk), .Q(mode_adj_654[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i2.GSR = "DISABLED";
    FD1P3IX SLO__i29 (.D(SLO[27]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i29.GSR = "DISABLED";
    FD1P3IX SLO__i30 (.D(SLO[28]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i30.GSR = "DISABLED";
    FD1P3IX SLO__i31 (.D(SLO[29]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i31.GSR = "DISABLED";
    CCU2D Cnt_NSL_1778_add_4_13 (.A0(Cnt_NSL[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21906), .S0(n53[11]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778_add_4_13.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1778_add_4_13.INIT1 = 16'h0000;
    defparam Cnt_NSL_1778_add_4_13.INJECT1_0 = "NO";
    defparam Cnt_NSL_1778_add_4_13.INJECT1_1 = "NO";
    FD1P3IX SLO__i32 (.D(SLO[30]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i32.GSR = "DISABLED";
    CCU2D Cnt_NSL_1778_add_4_11 (.A0(Cnt_NSL[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Cnt_NSL[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21905), .COUT(n21906), .S0(n53[9]), .S1(n53[10]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778_add_4_11.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1778_add_4_11.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1778_add_4_11.INJECT1_0 = "NO";
    defparam Cnt_NSL_1778_add_4_11.INJECT1_1 = "NO";
    FD1P3IX SLO__i33 (.D(SLO[31]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i33.GSR = "DISABLED";
    LUT4 i23949_4_lut (.A(NSL), .B(n30078), .C(n18522), .D(n30005), 
         .Z(NSL_N_4157)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C+(D))))) */ ;
    defparam i23949_4_lut.init = 16'h3b37;
    LUT4 i12769_2_lut_3_lut (.A(n18584), .B(n18522), .C(n153[1]), .Z(n199[1])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i12769_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_4_lut_adj_835 (.A(clk_enable_761), .B(EM_STOP), .C(n25721), 
         .D(n23916), .Z(clk_enable_1104)) /* synthesis lut_function=(A+!((C (D))+!B)) */ ;
    defparam i1_4_lut_adj_835.init = 16'haeee;
    CCU2D Cnt_NSL_1778_add_4_9 (.A0(Cnt_NSL[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Cnt_NSL[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21904), .COUT(n21905), .S0(n53[7]), .S1(n53[8]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778_add_4_9.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1778_add_4_9.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1778_add_4_9.INJECT1_0 = "NO";
    defparam Cnt_NSL_1778_add_4_9.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1778_add_4_7 (.A0(n93[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21903), .COUT(n21904), .S0(n53[5]), .S1(n53[6]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778_add_4_7.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1778_add_4_7.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1778_add_4_7.INJECT1_0 = "NO";
    defparam Cnt_NSL_1778_add_4_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_836 (.A(mode_adj_654[0]), .B(mode_adj_654[1]), .C(Cnt[4]), 
         .D(n4), .Z(n26363)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_836.init = 16'h8880;
    LUT4 i23892_1_lut_4_lut (.A(MA_Temp), .B(n18584), .C(n28326), .D(n30056), 
         .Z(n28586)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A (B+((D)+!C)))) */ ;
    defparam i23892_1_lut_4_lut.init = 16'h2212;
    CCU2D Cnt_NSL_1778_add_4_5 (.A0(n93[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21902), .COUT(n21903), .S0(n53[3]), .S1(n53[4]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778_add_4_5.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1778_add_4_5.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1778_add_4_5.INJECT1_0 = "NO";
    defparam Cnt_NSL_1778_add_4_5.INJECT1_1 = "NO";
    LUT4 i14080_2_lut_4_lut (.A(Cnt[1]), .B(n30131), .C(Cnt[0]), .D(Cnt[4]), 
         .Z(n18404)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam i14080_2_lut_4_lut.init = 16'hec00;
    LUT4 i14073_3_lut_4_lut (.A(n30177), .B(n30176), .C(resetn_c), .D(n18522), 
         .Z(clk_1MHz_enable_65)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i14073_3_lut_4_lut.init = 16'h70f0;
    CCU2D Cnt_NSL_1778_add_4_3 (.A0(n93[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21901), .COUT(n21902), .S0(n53[1]), .S1(n53[2]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778_add_4_3.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1778_add_4_3.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1778_add_4_3.INJECT1_0 = "NO";
    defparam Cnt_NSL_1778_add_4_3.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1778_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n30176), .B1(n30177), .C1(n93[0]), .D1(GND_net), 
          .COUT(n21901), .S1(n53[0]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1778_add_4_1.INIT0 = 16'hF000;
    defparam Cnt_NSL_1778_add_4_1.INIT1 = 16'h8787;
    defparam Cnt_NSL_1778_add_4_1.INJECT1_0 = "NO";
    defparam Cnt_NSL_1778_add_4_1.INJECT1_1 = "NO";
    LUT4 i23956_4_lut (.A(n25547), .B(n24169), .C(n18440), .D(n28402), 
         .Z(clk_enable_212)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i23956_4_lut.init = 16'hfff7;
    LUT4 mux_158_i36_3_lut (.A(SLO_buf[9]), .B(SLO_buf[3]), .C(n47), .Z(spi_data_out_r_39__N_4076[35])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i36_3_lut.init = 16'hcaca;
    LUT4 mux_158_i35_3_lut (.A(SLO_buf[8]), .B(SLO_buf[2]), .C(n47), .Z(spi_data_out_r_39__N_4076[34])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i35_3_lut.init = 16'hcaca;
    LUT4 mux_158_i34_3_lut (.A(SLO_buf[7]), .B(SLO_buf[1]), .C(n47), .Z(spi_data_out_r_39__N_4076[33])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i34_3_lut.init = 16'hcaca;
    LUT4 mux_158_i33_3_lut (.A(SLO_buf[6]), .B(SLO_buf[0]), .C(n47), .Z(spi_data_out_r_39__N_4076[32])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i33_3_lut.init = 16'hcaca;
    LUT4 mux_158_i16_3_lut (.A(SLO_buf[29]), .B(SLO_buf[19]), .C(n47), 
         .Z(spi_data_out_r_39__N_4076[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i16_3_lut.init = 16'hcaca;
    LUT4 mux_158_i15_3_lut (.A(SLO_buf[28]), .B(SLO_buf[18]), .C(n47), 
         .Z(spi_data_out_r_39__N_4076[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i15_3_lut.init = 16'hcaca;
    LUT4 mux_158_i14_3_lut (.A(SLO_buf[27]), .B(SLO_buf[17]), .C(n47), 
         .Z(spi_data_out_r_39__N_4076[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i14_3_lut.init = 16'hcaca;
    LUT4 mux_158_i13_3_lut (.A(SLO_buf[26]), .B(SLO_buf[16]), .C(n47), 
         .Z(spi_data_out_r_39__N_4076[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i13_3_lut.init = 16'hcaca;
    LUT4 mux_158_i12_3_lut (.A(SLO_buf[25]), .B(SLO_buf[15]), .C(n47), 
         .Z(spi_data_out_r_39__N_4076[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i12_3_lut.init = 16'hcaca;
    LUT4 mux_158_i11_3_lut (.A(SLO_buf[24]), .B(SLO_buf[14]), .C(n47), 
         .Z(spi_data_out_r_39__N_4076[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i11_3_lut.init = 16'hcaca;
    LUT4 mux_158_i10_3_lut (.A(SLO_buf[23]), .B(SLO_buf[13]), .C(n47), 
         .Z(spi_data_out_r_39__N_4076[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i10_3_lut.init = 16'hcaca;
    LUT4 mux_158_i9_3_lut (.A(SLO_buf[22]), .B(SLO_buf[12]), .C(n47), 
         .Z(spi_data_out_r_39__N_4076[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i9_3_lut.init = 16'hcaca;
    LUT4 mux_158_i8_3_lut (.A(SLO_buf[21]), .B(SLO_buf[11]), .C(n47), 
         .Z(spi_data_out_r_39__N_4076[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i8_3_lut.init = 16'hcaca;
    LUT4 mux_158_i7_3_lut (.A(SLO_buf[20]), .B(SLO_buf[10]), .C(n47), 
         .Z(spi_data_out_r_39__N_4076[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i7_3_lut.init = 16'hcaca;
    LUT4 mux_158_i6_3_lut (.A(SLO_buf[19]), .B(SLO_buf[9]), .C(n47), .Z(spi_data_out_r_39__N_4076[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i6_3_lut.init = 16'hcaca;
    LUT4 mux_158_i5_3_lut (.A(SLO_buf[18]), .B(SLO_buf[8]), .C(n47), .Z(spi_data_out_r_39__N_4076[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i5_3_lut.init = 16'hcaca;
    LUT4 mux_158_i4_3_lut (.A(SLO_buf[17]), .B(SLO_buf[7]), .C(n47), .Z(spi_data_out_r_39__N_4076[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i4_3_lut.init = 16'hcaca;
    LUT4 mux_158_i3_3_lut (.A(SLO_buf[16]), .B(SLO_buf[6]), .C(n47), .Z(spi_data_out_r_39__N_4076[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i3_3_lut.init = 16'hcaca;
    LUT4 mux_158_i2_3_lut (.A(SLO_buf[15]), .B(SLO_buf[5]), .C(n47), .Z(spi_data_out_r_39__N_4076[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i2_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_rep_599 (.A(n23916), .B(n28524), .C(n30045), .Z(n29999)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut_rep_599.init = 16'h2020;
    LUT4 i1_4_lut_adj_837 (.A(n28486), .B(n30045), .C(\spi_addr_r[4] ), 
         .D(\spi_addr_r[2] ), .Z(n27013)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_837.init = 16'h0400;
    LUT4 i1_2_lut_rep_772 (.A(\spi_addr_r[0] ), .B(\spi_cmd_r[0] ), .Z(n30172)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_772.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\spi_addr_r[0] ), .B(\spi_cmd_r[0] ), 
         .C(spi_data_valid_r), .D(\spi_addr_r[3] ), .Z(n25471)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2437_2_lut_rep_775 (.A(mode_adj_654[0]), .B(mode_adj_654[1]), 
         .Z(n30175)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2437_2_lut_rep_775.init = 16'h8888;
    LUT4 i2417_2_lut_rep_652_3_lut (.A(mode_adj_654[0]), .B(mode_adj_654[1]), 
         .C(mode_adj_654[2]), .Z(n30052)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i2417_2_lut_rep_652_3_lut.init = 16'hf8f8;
    LUT4 i1_3_lut_rep_776 (.A(Cnt_NSL[9]), .B(Cnt_NSL[8]), .C(Cnt_NSL[7]), 
         .Z(n30176)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_rep_776.init = 16'hfefe;
    LUT4 i1_2_lut_rep_678_4_lut (.A(Cnt_NSL[9]), .B(Cnt_NSL[8]), .C(Cnt_NSL[7]), 
         .D(n30177), .Z(n30078)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_rep_678_4_lut.init = 16'hfe00;
    LUT4 i1_2_lut_rep_777 (.A(Cnt_NSL[11]), .B(Cnt_NSL[10]), .Z(n30177)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i1_2_lut_rep_777.init = 16'h8888;
    LUT4 i23943_2_lut_rep_629_3_lut_4_lut (.A(Cnt_NSL[11]), .B(Cnt_NSL[10]), 
         .C(resetn_c), .D(n30176), .Z(clk_1MHz_enable_56)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i23943_2_lut_rep_629_3_lut_4_lut.init = 16'h8f0f;
    LUT4 i13290_2_lut_rep_790 (.A(Cnt[1]), .B(Cnt[4]), .Z(n30190)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13290_2_lut_rep_790.init = 16'h8888;
    LUT4 i1_2_lut_rep_605_3_lut_4_lut (.A(Cnt[1]), .B(Cnt[4]), .C(n30056), 
         .D(Cnt[5]), .Z(n30005)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_rep_605_3_lut_4_lut.init = 16'hfff7;
    LUT4 i23624_2_lut_3_lut (.A(Cnt[1]), .B(Cnt[4]), .C(Cnt[5]), .Z(n28326)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i23624_2_lut_3_lut.init = 16'h8080;
    LUT4 i12766_2_lut_3_lut (.A(n18584), .B(n18522), .C(n153[2]), .Z(n199[2])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i12766_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_607 (.A(n27013), .B(n23916), .Z(n30007)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_607.init = 16'h8888;
    LUT4 i24141_2_lut (.A(resetn_c), .B(n18440), .Z(clk_enable_242)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i24141_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_rep_594_3_lut (.A(n27013), .B(n23916), .C(n18440), .Z(n29994)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_594_3_lut.init = 16'h0808;
    FD1P3IX SLO__i34 (.D(SLO[32]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i34.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_799 (.A(\spi_addr_r[1] ), .B(\spi_cmd_r[2] ), .C(\spi_cmd_r[0] ), 
         .Z(n30199)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut_rep_799.init = 16'h1010;
    LUT4 i1_2_lut_4_lut_adj_838 (.A(\spi_addr_r[1] ), .B(\spi_cmd_r[2] ), 
         .C(\spi_cmd_r[0] ), .D(n25739), .Z(n25699)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_4_lut_adj_838.init = 16'h1000;
    LUT4 i1_2_lut_4_lut_adj_839 (.A(\spi_addr_r[1] ), .B(\spi_cmd_r[2] ), 
         .C(\spi_cmd_r[0] ), .D(n25941), .Z(n25943)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_4_lut_adj_839.init = 16'h1000;
    FD1P3IX SLO__i35 (.D(SLO[33]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i35.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_840 (.A(n23916), .B(n30109), .C(\spi_addr_r[1] ), 
         .D(n25793), .Z(n25801)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_840.init = 16'h0200;
    LUT4 i1_3_lut_adj_841 (.A(\spi_cmd_r[0] ), .B(\spi_addr_r[0] ), .C(resetn_c), 
         .Z(n25793)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_841.init = 16'h8080;
    LUT4 i1_3_lut_4_lut (.A(\spi_cmd_r[3] ), .B(n30044), .C(n26957), .D(n23916), 
         .Z(clk_enable_256)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut (.A(Cnt[5]), .B(n30056), .C(Cnt[1]), .Z(n4)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i23891_1_lut_2_lut_3_lut_4_lut (.A(Cnt[5]), .B(n30056), .C(MA_Temp), 
         .D(n30190), .Z(n28585)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam i23891_1_lut_2_lut_3_lut_4_lut.init = 16'he1f0;
    LUT4 i24039_2_lut_3_lut_4_lut (.A(resetn_c), .B(n30078), .C(n18522), 
         .D(n18584), .Z(clk_1MHz_enable_7)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (C (D)))) */ ;
    defparam i24039_2_lut_3_lut_4_lut.init = 16'h0ddd;
    LUT4 i23676_2_lut_rep_709 (.A(\spi_addr_r[3] ), .B(\spi_cmd_r[2] ), 
         .Z(n30109)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23676_2_lut_rep_709.init = 16'heeee;
    LUT4 i1_3_lut_rep_645_4_lut (.A(\spi_addr_r[3] ), .B(\spi_cmd_r[2] ), 
         .C(n30172), .D(\spi_addr_r[1] ), .Z(n30045)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_3_lut_rep_645_4_lut.init = 16'h0010;
    LUT4 i12757_2_lut_3_lut (.A(n18584), .B(n18522), .C(n153[6]), .Z(n199[6])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i12757_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_4_lut_adj_842 (.A(\spi_cmd_r[1] ), .B(\spi_cmd_r[4] ), .C(\spi_cmd_r[3] ), 
         .D(\spi_cmd_r[5] ), .Z(n18440)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_842.init = 16'hfffe;
    FD1P3AX NSL_484 (.D(NSL_N_4157), .SP(clk_1MHz_enable_65), .CK(clk_1MHz), 
            .Q(NSL)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam NSL_484.GSR = "DISABLED";
    FD1P3IX reset_r_491 (.D(reset_r_N_4129), .SP(clk_enable_1104), .CD(n30185), 
            .CK(clk), .Q(reset_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam reset_r_491.GSR = "DISABLED";
    FD1P3IX SLO__i36 (.D(SLO[34]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i36.GSR = "DISABLED";
    FD1P3IX SLO__i37 (.D(SLO[35]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i37.GSR = "DISABLED";
    CCU2D add_564_9 (.A0(Cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21917), 
          .S0(n153[7]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_9.INIT0 = 16'h5aaa;
    defparam add_564_9.INIT1 = 16'h0000;
    defparam add_564_9.INJECT1_0 = "NO";
    defparam add_564_9.INJECT1_1 = "NO";
    LUT4 i12750_2_lut_3_lut (.A(n18584), .B(n18522), .C(n153[7]), .Z(n199[7])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i12750_2_lut_3_lut.init = 16'h7070;
    FD1P3IX SLO__i38 (.D(SLO[36]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i38.GSR = "DISABLED";
    LUT4 i12761_2_lut_3_lut (.A(n18584), .B(n18522), .C(n153[5]), .Z(n199[5])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i12761_2_lut_3_lut.init = 16'h7070;
    FD1P3IX SLO__i39 (.D(SLO[37]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i39.GSR = "DISABLED";
    CCU2D add_564_7 (.A0(Cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21916), 
          .COUT(n21917), .S0(n153[5]), .S1(n153[6]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_7.INIT0 = 16'h5aaa;
    defparam add_564_7.INIT1 = 16'h5aaa;
    defparam add_564_7.INJECT1_0 = "NO";
    defparam add_564_7.INJECT1_1 = "NO";
    LUT4 i23953_2_lut_rep_729 (.A(MA_Temp), .B(clk_1MHz), .Z(n30129)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i23953_2_lut_rep_729.init = 16'h7777;
    LUT4 i12762_2_lut_3_lut (.A(n18584), .B(n18522), .C(n153[4]), .Z(n199[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i12762_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_663_3_lut (.A(MA_Temp), .B(clk_1MHz), .C(prev_MA), 
         .Z(n30063)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i1_2_lut_rep_663_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_730 (.A(Cnt[6]), .B(Cnt[7]), .Z(n30130)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam i1_2_lut_rep_730.init = 16'heeee;
    LUT4 i1_3_lut_rep_656_4_lut (.A(Cnt[6]), .B(Cnt[7]), .C(Cnt[0]), .D(n30131), 
         .Z(n30056)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam i1_3_lut_rep_656_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_731 (.A(Cnt[2]), .B(Cnt[3]), .Z(n30131)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam i1_2_lut_rep_731.init = 16'heeee;
    LUT4 i1_3_lut_rep_677_4_lut (.A(Cnt[2]), .B(Cnt[3]), .C(Cnt[0]), .D(Cnt[1]), 
         .Z(n30077)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam i1_3_lut_rep_677_4_lut.init = 16'hfeee;
    FD1P3IX SLO__i40 (.D(SLO[38]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i40.GSR = "DISABLED";
    FD1P3IX SLO__i41 (.D(SLO[39]), .SP(clk_enable_1132), .CD(n12235), 
            .CK(clk), .Q(SLO[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i41.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_734 (.A(mode_adj_654[1]), .B(mode_adj_654[0]), .Z(n30134)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_rep_734.init = 16'heeee;
    LUT4 i1_2_lut_rep_643_3_lut (.A(mode_adj_654[1]), .B(mode_adj_654[0]), 
         .C(mode_adj_654[2]), .Z(n30043)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_rep_643_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_618_3_lut_4_lut (.A(mode_adj_654[1]), .B(mode_adj_654[0]), 
         .C(mode_adj_653), .D(mode_adj_654[2]), .Z(n30018)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_rep_618_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2968_2_lut_3_lut_4_lut (.A(mode_adj_654[1]), .B(mode_adj_654[0]), 
         .C(pin_io_out_4), .D(mode_adj_654[2]), .Z(\pin_intrpt[2] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2968_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_2_lut_rep_658_3_lut (.A(mode_adj_654[1]), .B(mode_adj_654[0]), 
         .C(mode_adj_654[2]), .Z(n30058)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_rep_658_3_lut.init = 16'hefef;
    LUT4 i1_2_lut (.A(\quad_homing[0] ), .B(pin_io_out_4), .Z(n25869)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(74[8:17])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i12902_2_lut_3_lut (.A(n18584), .B(n18522), .C(n153[0]), .Z(n199[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i12902_2_lut_3_lut.init = 16'h7070;
    LUT4 i12763_2_lut_3_lut (.A(n18584), .B(n18522), .C(n153[3]), .Z(n199[3])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i12763_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_751 (.A(\spi_cmd_r[2] ), .B(\spi_cmd_r[0] ), .Z(n30151)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_rep_751.init = 16'h4444;
    LUT4 i1_3_lut_4_lut_adj_843 (.A(\spi_cmd_r[2] ), .B(\spi_cmd_r[0] ), 
         .C(\spi_addr_r[3] ), .D(n23916), .Z(n24169)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_3_lut_4_lut_adj_843.init = 16'h0400;
    
endmodule
//
// Verilog Description of module \quad_decoder(DEV_ID=3) 
//

module \quad_decoder(DEV_ID=3)  (n47, clk, n30185, \quad_b[3] , \spi_data_out_r_39__N_1639[0] , 
            \pin_intrpt[11] , \quad_a[3] , quad_homing, clk_enable_687, 
            \spi_data_r[0] , clk_enable_727, spi_data_out_r_39__N_1679, 
            spi_data_out_r_39__N_1868, n29990, \spi_data_out_r_39__N_1639[31] , 
            \spi_data_out_r_39__N_1639[30] , \spi_data_out_r_39__N_1639[29] , 
            \spi_data_out_r_39__N_1639[28] , \spi_data_out_r_39__N_1639[27] , 
            \spi_data_out_r_39__N_1639[26] , \spi_data_out_r_39__N_1639[25] , 
            \spi_data_out_r_39__N_1639[24] , \spi_data_out_r_39__N_1639[23] , 
            \spi_data_out_r_39__N_1639[22] , \spi_data_out_r_39__N_1639[21] , 
            \spi_data_out_r_39__N_1639[20] , \spi_data_out_r_39__N_1639[19] , 
            \spi_data_out_r_39__N_1639[18] , \spi_data_out_r_39__N_1639[17] , 
            \spi_data_out_r_39__N_1639[16] , \spi_data_out_r_39__N_1639[15] , 
            \spi_data_out_r_39__N_1639[14] , \spi_data_out_r_39__N_1639[13] , 
            \spi_data_out_r_39__N_1639[12] , \spi_data_out_r_39__N_1639[11] , 
            \spi_data_out_r_39__N_1639[10] , \spi_data_out_r_39__N_1639[9] , 
            \spi_data_out_r_39__N_1639[8] , \spi_data_out_r_39__N_1639[7] , 
            \spi_data_out_r_39__N_1639[6] , \spi_data_out_r_39__N_1639[5] , 
            \spi_data_out_r_39__N_1639[4] , \spi_data_out_r_39__N_1639[3] , 
            \spi_data_out_r_39__N_1639[2] , \spi_data_out_r_39__N_1639[1] , 
            n1, \spi_data_r[1] , \spi_data_r[2] , \spi_data_r[3] , \spi_data_r[4] , 
            \spi_data_r[5] , \spi_data_r[6] , \spi_data_r[7] , \spi_data_r[8] , 
            \spi_data_r[9] , \spi_data_r[10] , \spi_data_r[11] , \spi_data_r[12] , 
            \spi_data_r[13] , \spi_data_r[14] , \spi_data_r[15] , \spi_data_r[16] , 
            \spi_data_r[17] , \spi_data_r[18] , \spi_data_r[19] , \spi_data_r[20] , 
            \spi_data_r[21] , \spi_data_r[22] , \spi_data_r[23] , \spi_data_r[24] , 
            \spi_data_r[25] , \spi_data_r[26] , \spi_data_r[27] , \spi_data_r[28] , 
            \spi_data_r[29] , \spi_data_r[30] , \spi_data_r[31] , resetn_c, 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input n47;
    input clk;
    input n30185;
    input \quad_b[3] ;
    output \spi_data_out_r_39__N_1639[0] ;
    input \pin_intrpt[11] ;
    input \quad_a[3] ;
    output [1:0]quad_homing;
    input clk_enable_687;
    input \spi_data_r[0] ;
    input clk_enable_727;
    output spi_data_out_r_39__N_1679;
    input spi_data_out_r_39__N_1868;
    input n29990;
    output \spi_data_out_r_39__N_1639[31] ;
    output \spi_data_out_r_39__N_1639[30] ;
    output \spi_data_out_r_39__N_1639[29] ;
    output \spi_data_out_r_39__N_1639[28] ;
    output \spi_data_out_r_39__N_1639[27] ;
    output \spi_data_out_r_39__N_1639[26] ;
    output \spi_data_out_r_39__N_1639[25] ;
    output \spi_data_out_r_39__N_1639[24] ;
    output \spi_data_out_r_39__N_1639[23] ;
    output \spi_data_out_r_39__N_1639[22] ;
    output \spi_data_out_r_39__N_1639[21] ;
    output \spi_data_out_r_39__N_1639[20] ;
    output \spi_data_out_r_39__N_1639[19] ;
    output \spi_data_out_r_39__N_1639[18] ;
    output \spi_data_out_r_39__N_1639[17] ;
    output \spi_data_out_r_39__N_1639[16] ;
    output \spi_data_out_r_39__N_1639[15] ;
    output \spi_data_out_r_39__N_1639[14] ;
    output \spi_data_out_r_39__N_1639[13] ;
    output \spi_data_out_r_39__N_1639[12] ;
    output \spi_data_out_r_39__N_1639[11] ;
    output \spi_data_out_r_39__N_1639[10] ;
    output \spi_data_out_r_39__N_1639[9] ;
    output \spi_data_out_r_39__N_1639[8] ;
    output \spi_data_out_r_39__N_1639[7] ;
    output \spi_data_out_r_39__N_1639[6] ;
    output \spi_data_out_r_39__N_1639[5] ;
    output \spi_data_out_r_39__N_1639[4] ;
    output \spi_data_out_r_39__N_1639[3] ;
    output \spi_data_out_r_39__N_1639[2] ;
    output \spi_data_out_r_39__N_1639[1] ;
    input n1;
    input \spi_data_r[1] ;
    input \spi_data_r[2] ;
    input \spi_data_r[3] ;
    input \spi_data_r[4] ;
    input \spi_data_r[5] ;
    input \spi_data_r[6] ;
    input \spi_data_r[7] ;
    input \spi_data_r[8] ;
    input \spi_data_r[9] ;
    input \spi_data_r[10] ;
    input \spi_data_r[11] ;
    input \spi_data_r[12] ;
    input \spi_data_r[13] ;
    input \spi_data_r[14] ;
    input \spi_data_r[15] ;
    input \spi_data_r[16] ;
    input \spi_data_r[17] ;
    input \spi_data_r[18] ;
    input \spi_data_r[19] ;
    input \spi_data_r[20] ;
    input \spi_data_r[21] ;
    input \spi_data_r[22] ;
    input \spi_data_r[23] ;
    input \spi_data_r[24] ;
    input \spi_data_r[25] ;
    input \spi_data_r[26] ;
    input \spi_data_r[27] ;
    input \spi_data_r[28] ;
    input \spi_data_r[29] ;
    input \spi_data_r[30] ;
    input \spi_data_r[31] ;
    input resetn_c;
    input GND_net;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire \pin_intrpt[11]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[11] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    wire [31:0]quad_count;   // c:/s_links/sources/quad_decoder.v(43[29:39])
    wire [31:0]quad_buffer;   // c:/s_links/sources/quad_decoder.v(44[29:40])
    wire [39:0]spi_data_out_r_39__N_1788;
    
    wire clk_enable_453, n8533;
    wire [2:0]quad_b_delayed;   // c:/s_links/sources/quad_decoder.v(35[19:33])
    wire [2:0]quad_a_delayed;   // c:/s_links/sources/quad_decoder.v(34[20:34])
    wire [31:0]quad_set;   // c:/s_links/sources/quad_decoder.v(39[31:39])
    
    wire quad_set_valid, n9635, n9633, n9631, n9629, n9627, n9625, 
        n9623, n9621, n9619, n9617, n9615, n9613, n9611, n9609, 
        n9607, n9605, n9603, n9601, n9599, n9597, n9595, n9593, 
        n9591, n9589, n9587, n9585, n9583, n9581, n9579, n9577, 
        n9575;
    wire [31:0]n3996;
    
    wire n5705, n6, count_dir, n22059, n22058, n22057, n22056, 
        n22055, n22054, n22053, n22052, n22051, n22050, n22049, 
        n22048, n22047, n22046, n22045, n22044;
    
    LUT4 mux_425_i7_3_lut (.A(quad_count[6]), .B(quad_buffer[6]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i7_3_lut.init = 16'hcaca;
    FD1P3AX quad_count_i0_i0 (.D(n8533), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i0.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i0 (.D(\quad_b[3] ), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(spi_data_out_r_39__N_1788[0]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX quad_buffer_i0 (.D(quad_count[0]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i0.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i0 (.D(\quad_a[3] ), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i0.GSR = "DISABLED";
    FD1P3IX quad_homing__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_687), .CD(n30185), 
            .CK(clk), .Q(quad_homing[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(62[8] 69[4])
    defparam quad_homing__i0.GSR = "DISABLED";
    FD1P3IX quad_set__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i0.GSR = "DISABLED";
    LUT4 mux_425_i6_3_lut (.A(quad_count[5]), .B(quad_buffer[5]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i6_3_lut.init = 16'hcaca;
    LUT4 mux_425_i5_3_lut (.A(quad_count[4]), .B(quad_buffer[4]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i5_3_lut.init = 16'hcaca;
    LUT4 mux_425_i4_3_lut (.A(quad_count[3]), .B(quad_buffer[3]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i4_3_lut.init = 16'hcaca;
    LUT4 mux_425_i3_3_lut (.A(quad_count[2]), .B(quad_buffer[2]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i3_3_lut.init = 16'hcaca;
    LUT4 mux_425_i2_3_lut (.A(quad_count[1]), .B(quad_buffer[1]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i2_3_lut.init = 16'hcaca;
    FD1S3IX i39_391 (.D(spi_data_out_r_39__N_1868), .CK(clk), .CD(n30185), 
            .Q(spi_data_out_r_39__N_1679)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam i39_391.GSR = "DISABLED";
    FD1S3IX quad_set_valid_388 (.D(n29990), .CK(clk), .CD(n30185), .Q(quad_set_valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set_valid_388.GSR = "DISABLED";
    FD1S3AX quad_buffer_i31 (.D(quad_count[31]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i31.GSR = "DISABLED";
    FD1S3AX quad_buffer_i30 (.D(quad_count[30]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i30.GSR = "DISABLED";
    FD1S3AX quad_buffer_i29 (.D(quad_count[29]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i29.GSR = "DISABLED";
    FD1S3AX quad_buffer_i28 (.D(quad_count[28]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i28.GSR = "DISABLED";
    FD1S3AX quad_buffer_i27 (.D(quad_count[27]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i27.GSR = "DISABLED";
    FD1S3AX quad_buffer_i26 (.D(quad_count[26]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i26.GSR = "DISABLED";
    FD1S3AX quad_buffer_i25 (.D(quad_count[25]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i25.GSR = "DISABLED";
    FD1S3AX quad_buffer_i24 (.D(quad_count[24]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i24.GSR = "DISABLED";
    FD1S3AX quad_buffer_i23 (.D(quad_count[23]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i23.GSR = "DISABLED";
    FD1S3AX quad_buffer_i22 (.D(quad_count[22]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i22.GSR = "DISABLED";
    FD1S3AX quad_buffer_i21 (.D(quad_count[21]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i21.GSR = "DISABLED";
    FD1S3AX quad_buffer_i20 (.D(quad_count[20]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i20.GSR = "DISABLED";
    FD1S3AX quad_buffer_i19 (.D(quad_count[19]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i19.GSR = "DISABLED";
    FD1S3AX quad_buffer_i18 (.D(quad_count[18]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i18.GSR = "DISABLED";
    FD1S3AX quad_buffer_i17 (.D(quad_count[17]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i17.GSR = "DISABLED";
    FD1S3AX quad_buffer_i16 (.D(quad_count[16]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i16.GSR = "DISABLED";
    FD1S3AX quad_buffer_i15 (.D(quad_count[15]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i15.GSR = "DISABLED";
    FD1S3AX quad_buffer_i14 (.D(quad_count[14]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i14.GSR = "DISABLED";
    FD1S3AX quad_buffer_i13 (.D(quad_count[13]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i13.GSR = "DISABLED";
    FD1S3AX quad_buffer_i12 (.D(quad_count[12]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i12.GSR = "DISABLED";
    FD1S3AX quad_buffer_i11 (.D(quad_count[11]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i11.GSR = "DISABLED";
    FD1S3AX quad_buffer_i10 (.D(quad_count[10]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i10.GSR = "DISABLED";
    FD1S3AX quad_buffer_i9 (.D(quad_count[9]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i9.GSR = "DISABLED";
    FD1S3AX quad_buffer_i8 (.D(quad_count[8]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i8.GSR = "DISABLED";
    FD1S3AX quad_buffer_i7 (.D(quad_count[7]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i7.GSR = "DISABLED";
    FD1S3AX quad_buffer_i6 (.D(quad_count[6]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i6.GSR = "DISABLED";
    FD1S3AX quad_buffer_i5 (.D(quad_count[5]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i5.GSR = "DISABLED";
    FD1S3AX quad_buffer_i4 (.D(quad_count[4]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i4.GSR = "DISABLED";
    FD1S3AX quad_buffer_i3 (.D(quad_count[3]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i3.GSR = "DISABLED";
    FD1S3AX quad_buffer_i2 (.D(quad_count[2]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i2.GSR = "DISABLED";
    FD1S3AX quad_buffer_i1 (.D(quad_count[1]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(spi_data_out_r_39__N_1788[31]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i31 (.D(spi_data_out_r_39__N_1788[30]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i30 (.D(spi_data_out_r_39__N_1788[29]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i29 (.D(spi_data_out_r_39__N_1788[28]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i28 (.D(spi_data_out_r_39__N_1788[27]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i27 (.D(spi_data_out_r_39__N_1788[26]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i26 (.D(spi_data_out_r_39__N_1788[25]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i25 (.D(spi_data_out_r_39__N_1788[24]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i24 (.D(spi_data_out_r_39__N_1788[23]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i23 (.D(spi_data_out_r_39__N_1788[22]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i22 (.D(spi_data_out_r_39__N_1788[21]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i21 (.D(spi_data_out_r_39__N_1788[20]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i20 (.D(spi_data_out_r_39__N_1788[19]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i19 (.D(spi_data_out_r_39__N_1788[18]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i18 (.D(spi_data_out_r_39__N_1788[17]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i17 (.D(spi_data_out_r_39__N_1788[16]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i16 (.D(spi_data_out_r_39__N_1788[15]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(spi_data_out_r_39__N_1788[14]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(spi_data_out_r_39__N_1788[13]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(spi_data_out_r_39__N_1788[12]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(spi_data_out_r_39__N_1788[11]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(spi_data_out_r_39__N_1788[10]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(spi_data_out_r_39__N_1788[9]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(spi_data_out_r_39__N_1788[8]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(spi_data_out_r_39__N_1788[7]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(spi_data_out_r_39__N_1788[6]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(spi_data_out_r_39__N_1788[5]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(spi_data_out_r_39__N_1788[4]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(spi_data_out_r_39__N_1788[3]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(spi_data_out_r_39__N_1788[2]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(spi_data_out_r_39__N_1788[1]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1639[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i2 (.D(quad_b_delayed[1]), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i2.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i1 (.D(quad_b_delayed[0]), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i1.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i31 (.D(n9635), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i31.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i30 (.D(n9633), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i30.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i29 (.D(n9631), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i29.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i28 (.D(n9629), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i28.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i27 (.D(n9627), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i27.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i26 (.D(n9625), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i26.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i25 (.D(n9623), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i25.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i24 (.D(n9621), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i24.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i23 (.D(n9619), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i23.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i22 (.D(n9617), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i22.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i21 (.D(n9615), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i21.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i20 (.D(n9613), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i20.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i19 (.D(n9611), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i19.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i18 (.D(n9609), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i18.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i17 (.D(n9607), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i17.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i16 (.D(n9605), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i16.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i15 (.D(n9603), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i15.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i14 (.D(n9601), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i14.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i13 (.D(n9599), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i13.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i12 (.D(n9597), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i12.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i11 (.D(n9595), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i11.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i10 (.D(n9593), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i10.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i9 (.D(n9591), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i9.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i8 (.D(n9589), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i8.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i7 (.D(n9587), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i7.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i6 (.D(n9585), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i6.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i5 (.D(n9583), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i5.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i4 (.D(n9581), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i4.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i3 (.D(n9579), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i3.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i2 (.D(n9577), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i1 (.D(n9575), .SP(clk_enable_453), .CK(clk), 
            .Q(quad_count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i1.GSR = "DISABLED";
    LUT4 i5297_4_lut (.A(n3996[24]), .B(quad_set[24]), .C(n5705), .D(n1), 
         .Z(n9621)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5297_4_lut.init = 16'hc0ca;
    LUT4 i5295_4_lut (.A(n3996[23]), .B(quad_set[23]), .C(n5705), .D(n1), 
         .Z(n9619)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5295_4_lut.init = 16'hc0ca;
    LUT4 i5293_4_lut (.A(n3996[22]), .B(quad_set[22]), .C(n5705), .D(n1), 
         .Z(n9617)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5293_4_lut.init = 16'hc0ca;
    LUT4 i5291_4_lut (.A(n3996[21]), .B(quad_set[21]), .C(n5705), .D(n1), 
         .Z(n9615)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5291_4_lut.init = 16'hc0ca;
    LUT4 i5289_4_lut (.A(n3996[20]), .B(quad_set[20]), .C(n5705), .D(n1), 
         .Z(n9613)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5289_4_lut.init = 16'hc0ca;
    LUT4 i5287_4_lut (.A(n3996[19]), .B(quad_set[19]), .C(n5705), .D(n1), 
         .Z(n9611)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5287_4_lut.init = 16'hc0ca;
    LUT4 i5285_4_lut (.A(n3996[18]), .B(quad_set[18]), .C(n5705), .D(n1), 
         .Z(n9609)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5285_4_lut.init = 16'hc0ca;
    LUT4 i5283_4_lut (.A(n3996[17]), .B(quad_set[17]), .C(n5705), .D(n1), 
         .Z(n9607)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5283_4_lut.init = 16'hc0ca;
    LUT4 i5281_4_lut (.A(n3996[16]), .B(quad_set[16]), .C(n5705), .D(n1), 
         .Z(n9605)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5281_4_lut.init = 16'hc0ca;
    LUT4 i5279_4_lut (.A(n3996[15]), .B(quad_set[15]), .C(n5705), .D(n1), 
         .Z(n9603)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5279_4_lut.init = 16'hc0ca;
    LUT4 i5277_4_lut (.A(n3996[14]), .B(quad_set[14]), .C(n5705), .D(n1), 
         .Z(n9601)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5277_4_lut.init = 16'hc0ca;
    LUT4 i5275_4_lut (.A(n3996[13]), .B(quad_set[13]), .C(n5705), .D(n1), 
         .Z(n9599)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5275_4_lut.init = 16'hc0ca;
    LUT4 i5273_4_lut (.A(n3996[12]), .B(quad_set[12]), .C(n5705), .D(n1), 
         .Z(n9597)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5273_4_lut.init = 16'hc0ca;
    LUT4 i5271_4_lut (.A(n3996[11]), .B(quad_set[11]), .C(n5705), .D(n1), 
         .Z(n9595)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5271_4_lut.init = 16'hc0ca;
    LUT4 i5269_4_lut (.A(n3996[10]), .B(quad_set[10]), .C(n5705), .D(n1), 
         .Z(n9593)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5269_4_lut.init = 16'hc0ca;
    LUT4 i5267_4_lut (.A(n3996[9]), .B(quad_set[9]), .C(n5705), .D(n1), 
         .Z(n9591)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5267_4_lut.init = 16'hc0ca;
    LUT4 i5265_4_lut (.A(n3996[8]), .B(quad_set[8]), .C(n5705), .D(n1), 
         .Z(n9589)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5265_4_lut.init = 16'hc0ca;
    LUT4 i5263_4_lut (.A(n3996[7]), .B(quad_set[7]), .C(n5705), .D(n1), 
         .Z(n9587)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5263_4_lut.init = 16'hc0ca;
    LUT4 i5261_4_lut (.A(n3996[6]), .B(quad_set[6]), .C(n5705), .D(n1), 
         .Z(n9585)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5261_4_lut.init = 16'hc0ca;
    LUT4 i5259_4_lut (.A(n3996[5]), .B(quad_set[5]), .C(n5705), .D(n1), 
         .Z(n9583)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5259_4_lut.init = 16'hc0ca;
    LUT4 i5257_4_lut (.A(n3996[4]), .B(quad_set[4]), .C(n5705), .D(n1), 
         .Z(n9581)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5257_4_lut.init = 16'hc0ca;
    LUT4 i5255_4_lut (.A(n3996[3]), .B(quad_set[3]), .C(n5705), .D(n1), 
         .Z(n9579)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5255_4_lut.init = 16'hc0ca;
    LUT4 i5253_4_lut (.A(n3996[2]), .B(quad_set[2]), .C(n5705), .D(n1), 
         .Z(n9577)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5253_4_lut.init = 16'hc0ca;
    LUT4 i5251_4_lut (.A(n3996[1]), .B(quad_set[1]), .C(n5705), .D(n1), 
         .Z(n9575)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5251_4_lut.init = 16'hc0ca;
    LUT4 i2_2_lut (.A(quad_b_delayed[1]), .B(quad_a_delayed[2]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(96[19:96])
    defparam i2_2_lut.init = 16'h6666;
    LUT4 i1_2_lut (.A(quad_a_delayed[1]), .B(quad_b_delayed[2]), .Z(count_dir)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(96[19:96])
    defparam i1_2_lut.init = 16'h6666;
    FD1S3IX quad_a_delayed__i1 (.D(quad_a_delayed[0]), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i1.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i2 (.D(quad_a_delayed[1]), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i2.GSR = "DISABLED";
    FD1P3IX quad_homing__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_687), .CD(n30185), 
            .CK(clk), .Q(quad_homing[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(62[8] 69[4])
    defparam quad_homing__i1.GSR = "DISABLED";
    FD1P3IX quad_set__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i1.GSR = "DISABLED";
    FD1P3IX quad_set__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i2.GSR = "DISABLED";
    FD1P3IX quad_set__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i3.GSR = "DISABLED";
    FD1P3IX quad_set__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i4.GSR = "DISABLED";
    FD1P3IX quad_set__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i5.GSR = "DISABLED";
    FD1P3IX quad_set__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i6.GSR = "DISABLED";
    FD1P3IX quad_set__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i7.GSR = "DISABLED";
    FD1P3IX quad_set__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i8.GSR = "DISABLED";
    FD1P3IX quad_set__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i9.GSR = "DISABLED";
    FD1P3IX quad_set__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i10.GSR = "DISABLED";
    FD1P3IX quad_set__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i11.GSR = "DISABLED";
    FD1P3IX quad_set__i12 (.D(\spi_data_r[12] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i12.GSR = "DISABLED";
    FD1P3IX quad_set__i13 (.D(\spi_data_r[13] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i13.GSR = "DISABLED";
    FD1P3IX quad_set__i14 (.D(\spi_data_r[14] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i14.GSR = "DISABLED";
    FD1P3IX quad_set__i15 (.D(\spi_data_r[15] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i15.GSR = "DISABLED";
    FD1P3IX quad_set__i16 (.D(\spi_data_r[16] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i16.GSR = "DISABLED";
    FD1P3IX quad_set__i17 (.D(\spi_data_r[17] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i17.GSR = "DISABLED";
    FD1P3IX quad_set__i18 (.D(\spi_data_r[18] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i18.GSR = "DISABLED";
    FD1P3IX quad_set__i19 (.D(\spi_data_r[19] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i19.GSR = "DISABLED";
    FD1P3IX quad_set__i20 (.D(\spi_data_r[20] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i20.GSR = "DISABLED";
    FD1P3IX quad_set__i21 (.D(\spi_data_r[21] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i21.GSR = "DISABLED";
    FD1P3IX quad_set__i22 (.D(\spi_data_r[22] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i22.GSR = "DISABLED";
    FD1P3IX quad_set__i23 (.D(\spi_data_r[23] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i23.GSR = "DISABLED";
    FD1P3IX quad_set__i24 (.D(\spi_data_r[24] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i24.GSR = "DISABLED";
    FD1P3IX quad_set__i25 (.D(\spi_data_r[25] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i25.GSR = "DISABLED";
    FD1P3IX quad_set__i26 (.D(\spi_data_r[26] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i26.GSR = "DISABLED";
    FD1P3IX quad_set__i27 (.D(\spi_data_r[27] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i27.GSR = "DISABLED";
    FD1P3IX quad_set__i28 (.D(\spi_data_r[28] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i28.GSR = "DISABLED";
    FD1P3IX quad_set__i29 (.D(\spi_data_r[29] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i29.GSR = "DISABLED";
    FD1P3IX quad_set__i30 (.D(\spi_data_r[30] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i30.GSR = "DISABLED";
    FD1P3IX quad_set__i31 (.D(\spi_data_r[31] ), .SP(clk_enable_727), .CD(n30185), 
            .CK(clk), .Q(quad_set[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i31.GSR = "DISABLED";
    LUT4 i5299_4_lut (.A(n3996[25]), .B(quad_set[25]), .C(n5705), .D(n1), 
         .Z(n9623)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5299_4_lut.init = 16'hc0ca;
    LUT4 i24193_2_lut (.A(resetn_c), .B(quad_homing[1]), .Z(clk_enable_453)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i24193_2_lut.init = 16'h7777;
    LUT4 i4209_4_lut (.A(n3996[0]), .B(quad_set[0]), .C(n5705), .D(n1), 
         .Z(n8533)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4209_4_lut.init = 16'hc0ca;
    LUT4 i1_4_lut (.A(quad_homing[0]), .B(quad_homing[1]), .C(quad_set_valid), 
         .D(resetn_c), .Z(n5705)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut.init = 16'h1000;
    CCU2D add_1373_33 (.A0(quad_count[30]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[31]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22059), .S0(n3996[30]), .S1(n3996[31]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_33.INIT0 = 16'h5569;
    defparam add_1373_33.INIT1 = 16'h5569;
    defparam add_1373_33.INJECT1_0 = "NO";
    defparam add_1373_33.INJECT1_1 = "NO";
    CCU2D add_1373_31 (.A0(quad_count[28]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[29]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22058), .COUT(n22059), .S0(n3996[28]), .S1(n3996[29]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_31.INIT0 = 16'h5569;
    defparam add_1373_31.INIT1 = 16'h5569;
    defparam add_1373_31.INJECT1_0 = "NO";
    defparam add_1373_31.INJECT1_1 = "NO";
    CCU2D add_1373_29 (.A0(quad_count[26]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[27]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22057), .COUT(n22058), .S0(n3996[26]), .S1(n3996[27]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_29.INIT0 = 16'h5569;
    defparam add_1373_29.INIT1 = 16'h5569;
    defparam add_1373_29.INJECT1_0 = "NO";
    defparam add_1373_29.INJECT1_1 = "NO";
    CCU2D add_1373_27 (.A0(quad_count[24]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[25]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22056), .COUT(n22057), .S0(n3996[24]), .S1(n3996[25]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_27.INIT0 = 16'h5569;
    defparam add_1373_27.INIT1 = 16'h5569;
    defparam add_1373_27.INJECT1_0 = "NO";
    defparam add_1373_27.INJECT1_1 = "NO";
    CCU2D add_1373_25 (.A0(quad_count[22]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[23]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22055), .COUT(n22056), .S0(n3996[22]), .S1(n3996[23]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_25.INIT0 = 16'h5569;
    defparam add_1373_25.INIT1 = 16'h5569;
    defparam add_1373_25.INJECT1_0 = "NO";
    defparam add_1373_25.INJECT1_1 = "NO";
    CCU2D add_1373_23 (.A0(quad_count[20]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[21]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22054), .COUT(n22055), .S0(n3996[20]), .S1(n3996[21]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_23.INIT0 = 16'h5569;
    defparam add_1373_23.INIT1 = 16'h5569;
    defparam add_1373_23.INJECT1_0 = "NO";
    defparam add_1373_23.INJECT1_1 = "NO";
    CCU2D add_1373_21 (.A0(quad_count[18]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[19]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22053), .COUT(n22054), .S0(n3996[18]), .S1(n3996[19]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_21.INIT0 = 16'h5569;
    defparam add_1373_21.INIT1 = 16'h5569;
    defparam add_1373_21.INJECT1_0 = "NO";
    defparam add_1373_21.INJECT1_1 = "NO";
    CCU2D add_1373_19 (.A0(quad_count[16]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[17]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22052), .COUT(n22053), .S0(n3996[16]), .S1(n3996[17]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_19.INIT0 = 16'h5569;
    defparam add_1373_19.INIT1 = 16'h5569;
    defparam add_1373_19.INJECT1_0 = "NO";
    defparam add_1373_19.INJECT1_1 = "NO";
    CCU2D add_1373_17 (.A0(quad_count[14]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[15]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22051), .COUT(n22052), .S0(n3996[14]), .S1(n3996[15]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_17.INIT0 = 16'h5569;
    defparam add_1373_17.INIT1 = 16'h5569;
    defparam add_1373_17.INJECT1_0 = "NO";
    defparam add_1373_17.INJECT1_1 = "NO";
    CCU2D add_1373_15 (.A0(quad_count[12]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[13]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22050), .COUT(n22051), .S0(n3996[12]), .S1(n3996[13]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_15.INIT0 = 16'h5569;
    defparam add_1373_15.INIT1 = 16'h5569;
    defparam add_1373_15.INJECT1_0 = "NO";
    defparam add_1373_15.INJECT1_1 = "NO";
    CCU2D add_1373_13 (.A0(quad_count[10]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[11]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22049), .COUT(n22050), .S0(n3996[10]), .S1(n3996[11]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_13.INIT0 = 16'h5569;
    defparam add_1373_13.INIT1 = 16'h5569;
    defparam add_1373_13.INJECT1_0 = "NO";
    defparam add_1373_13.INJECT1_1 = "NO";
    CCU2D add_1373_11 (.A0(quad_count[8]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[9]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22048), .COUT(n22049), .S0(n3996[8]), .S1(n3996[9]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_11.INIT0 = 16'h5569;
    defparam add_1373_11.INIT1 = 16'h5569;
    defparam add_1373_11.INJECT1_0 = "NO";
    defparam add_1373_11.INJECT1_1 = "NO";
    CCU2D add_1373_9 (.A0(quad_count[6]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[7]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22047), .COUT(n22048), .S0(n3996[6]), .S1(n3996[7]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_9.INIT0 = 16'h5569;
    defparam add_1373_9.INIT1 = 16'h5569;
    defparam add_1373_9.INJECT1_0 = "NO";
    defparam add_1373_9.INJECT1_1 = "NO";
    CCU2D add_1373_7 (.A0(quad_count[4]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[5]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22046), .COUT(n22047), .S0(n3996[4]), .S1(n3996[5]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_7.INIT0 = 16'h5569;
    defparam add_1373_7.INIT1 = 16'h5569;
    defparam add_1373_7.INJECT1_0 = "NO";
    defparam add_1373_7.INJECT1_1 = "NO";
    CCU2D add_1373_5 (.A0(quad_count[2]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[3]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22045), .COUT(n22046), .S0(n3996[2]), .S1(n3996[3]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_5.INIT0 = 16'h5569;
    defparam add_1373_5.INIT1 = 16'h5569;
    defparam add_1373_5.INJECT1_0 = "NO";
    defparam add_1373_5.INJECT1_1 = "NO";
    CCU2D add_1373_3 (.A0(quad_count[0]), .B0(count_dir), .C0(n6), .D0(count_dir), 
          .A1(quad_count[1]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22044), .COUT(n22045), .S0(n3996[0]), .S1(n3996[1]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_3.INIT0 = 16'h5665;
    defparam add_1373_3.INIT1 = 16'h5569;
    defparam add_1373_3.INJECT1_0 = "NO";
    defparam add_1373_3.INJECT1_1 = "NO";
    CCU2D add_1373_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quad_a_delayed[2]), .B1(quad_b_delayed[1]), .C1(quad_b_delayed[2]), 
          .D1(quad_a_delayed[1]), .COUT(n22044));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1373_1.INIT0 = 16'hF000;
    defparam add_1373_1.INIT1 = 16'h0990;
    defparam add_1373_1.INJECT1_0 = "NO";
    defparam add_1373_1.INJECT1_1 = "NO";
    LUT4 mux_425_i1_3_lut (.A(quad_count[0]), .B(quad_buffer[0]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i1_3_lut.init = 16'hcaca;
    LUT4 mux_425_i32_3_lut (.A(quad_count[31]), .B(quad_buffer[31]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i32_3_lut.init = 16'hcaca;
    LUT4 mux_425_i31_3_lut (.A(quad_count[30]), .B(quad_buffer[30]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i31_3_lut.init = 16'hcaca;
    LUT4 mux_425_i30_3_lut (.A(quad_count[29]), .B(quad_buffer[29]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i30_3_lut.init = 16'hcaca;
    LUT4 mux_425_i29_3_lut (.A(quad_count[28]), .B(quad_buffer[28]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i29_3_lut.init = 16'hcaca;
    LUT4 mux_425_i28_3_lut (.A(quad_count[27]), .B(quad_buffer[27]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i28_3_lut.init = 16'hcaca;
    LUT4 mux_425_i27_3_lut (.A(quad_count[26]), .B(quad_buffer[26]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i27_3_lut.init = 16'hcaca;
    LUT4 mux_425_i26_3_lut (.A(quad_count[25]), .B(quad_buffer[25]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i26_3_lut.init = 16'hcaca;
    LUT4 mux_425_i25_3_lut (.A(quad_count[24]), .B(quad_buffer[24]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i25_3_lut.init = 16'hcaca;
    LUT4 mux_425_i24_3_lut (.A(quad_count[23]), .B(quad_buffer[23]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i24_3_lut.init = 16'hcaca;
    LUT4 mux_425_i23_3_lut (.A(quad_count[22]), .B(quad_buffer[22]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i23_3_lut.init = 16'hcaca;
    LUT4 mux_425_i22_3_lut (.A(quad_count[21]), .B(quad_buffer[21]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i22_3_lut.init = 16'hcaca;
    LUT4 mux_425_i21_3_lut (.A(quad_count[20]), .B(quad_buffer[20]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i21_3_lut.init = 16'hcaca;
    LUT4 mux_425_i20_3_lut (.A(quad_count[19]), .B(quad_buffer[19]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i20_3_lut.init = 16'hcaca;
    LUT4 mux_425_i19_3_lut (.A(quad_count[18]), .B(quad_buffer[18]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i19_3_lut.init = 16'hcaca;
    LUT4 mux_425_i18_3_lut (.A(quad_count[17]), .B(quad_buffer[17]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i18_3_lut.init = 16'hcaca;
    LUT4 mux_425_i17_3_lut (.A(quad_count[16]), .B(quad_buffer[16]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i17_3_lut.init = 16'hcaca;
    LUT4 mux_425_i16_3_lut (.A(quad_count[15]), .B(quad_buffer[15]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i16_3_lut.init = 16'hcaca;
    LUT4 mux_425_i15_3_lut (.A(quad_count[14]), .B(quad_buffer[14]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i15_3_lut.init = 16'hcaca;
    LUT4 mux_425_i14_3_lut (.A(quad_count[13]), .B(quad_buffer[13]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i14_3_lut.init = 16'hcaca;
    LUT4 mux_425_i13_3_lut (.A(quad_count[12]), .B(quad_buffer[12]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i13_3_lut.init = 16'hcaca;
    LUT4 mux_425_i12_3_lut (.A(quad_count[11]), .B(quad_buffer[11]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i12_3_lut.init = 16'hcaca;
    LUT4 mux_425_i11_3_lut (.A(quad_count[10]), .B(quad_buffer[10]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i11_3_lut.init = 16'hcaca;
    LUT4 mux_425_i9_3_lut (.A(quad_count[8]), .B(quad_buffer[8]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i9_3_lut.init = 16'hcaca;
    LUT4 mux_425_i8_3_lut (.A(quad_count[7]), .B(quad_buffer[7]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i8_3_lut.init = 16'hcaca;
    LUT4 mux_425_i10_3_lut (.A(quad_count[9]), .B(quad_buffer[9]), .C(n47), 
         .Z(spi_data_out_r_39__N_1788[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(77[7] 80[28])
    defparam mux_425_i10_3_lut.init = 16'hcaca;
    LUT4 i5311_4_lut (.A(n3996[31]), .B(quad_set[31]), .C(n5705), .D(n1), 
         .Z(n9635)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5311_4_lut.init = 16'hc0ca;
    LUT4 i5309_4_lut (.A(n3996[30]), .B(quad_set[30]), .C(n5705), .D(n1), 
         .Z(n9633)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5309_4_lut.init = 16'hc0ca;
    LUT4 i5307_4_lut (.A(n3996[29]), .B(quad_set[29]), .C(n5705), .D(n1), 
         .Z(n9631)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5307_4_lut.init = 16'hc0ca;
    LUT4 i5305_4_lut (.A(n3996[28]), .B(quad_set[28]), .C(n5705), .D(n1), 
         .Z(n9629)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5305_4_lut.init = 16'hc0ca;
    LUT4 i5303_4_lut (.A(n3996[27]), .B(quad_set[27]), .C(n5705), .D(n1), 
         .Z(n9627)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5303_4_lut.init = 16'hc0ca;
    LUT4 i5301_4_lut (.A(n3996[26]), .B(quad_set[26]), .C(n5705), .D(n1), 
         .Z(n9625)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5301_4_lut.init = 16'hc0ca;
    
endmodule
//
// Verilog Description of module \stepper(DEV_ID=3,UART_ADDRESS_WIDTH=4) 
//

module \stepper(DEV_ID=3,UART_ADDRESS_WIDTH=4)  (clk, GND_net, reset_r, 
            clk_enable_28, n30185, n29995, clk_1MHz, clk_enable_178, 
            \spi_data_r[0] , n30188, spi_data_out_r_39__N_4854, \spi_data_out_r_39__N_5105[0] , 
            resetn_c, \SLO_buf[0] , \spi_data_r[2] , \spi_data_r[1] , 
            spi_data_out_r_39__N_4894, spi_data_out_r_39__N_5191, digital_output_r, 
            clk_enable_254, n28554, pin_io_c_38, \spi_data_out_r_39__N_5105[1] , 
            \spi_data_out_r_39__N_5105[2] , \spi_data_out_r_39__N_5105[3] , 
            \spi_data_out_r_39__N_5105[4] , \spi_data_out_r_39__N_5105[5] , 
            \spi_data_out_r_39__N_5105[6] , \spi_data_out_r_39__N_5105[7] , 
            \spi_data_out_r_39__N_5105[8] , \spi_data_out_r_39__N_5105[9] , 
            \spi_data_out_r_39__N_5105[10] , \spi_data_out_r_39__N_5105[11] , 
            \spi_data_out_r_39__N_5105[12] , \spi_data_out_r_39__N_5105[13] , 
            \spi_data_out_r_39__N_5105[14] , \spi_data_out_r_39__N_5105[15] , 
            n29991, \spi_data_out_r_39__N_5105[32] , \spi_data_out_r_39__N_5105[33] , 
            \spi_data_out_r_39__N_5105[34] , \spi_data_out_r_39__N_5105[35] , 
            \SLO_buf[10] , \SLO_buf[11] , \SLO_buf[12] , \SLO_buf[13] , 
            \SLO_buf[1] , \SLO_buf[2] , \SLO_buf[3] , \SLO_buf[4] , 
            \SLO_buf[5] , \SLO_buf[6] , \SLO_buf[7] , \SLO_buf[8] , 
            \SLO_buf[9] , \SLO_buf[14] , \SLO_buf[15] , \SLO_buf[16] , 
            \SLO_buf[17] , \SLO_buf[18] , \SLO_buf[19] , \SLO_buf[20] , 
            \SLO_buf[21] , \SLO_buf[22] , \SLO_buf[23] , \SLO_buf[24] , 
            \SLO_buf[25] , \SLO_buf[26] , \SLO_buf[27] , \SLO_buf[28] , 
            \SLO_buf[29] , NSL, \quad_homing[0] , pin_io_c_34, n25873, 
            mode, \cs_decoded[6] , n7170, n30082, n7166, n30091, 
            pin_io_out_35, n29943, pin_io_c_33, \pin_intrpt[10] , pin_io_c_32, 
            \pin_intrpt[9] , \pin_intrpt[11] , n7269, UC_TXD0_c, OW_ID_N_5147, 
            n30050, ENC_O_N_5155, OW_ID_N_5153, \quad_a[3] , pin_io_out_39, 
            \quad_b[3] , \uart_slot_en[1] , \uart_slot_en[0] , n10696, 
            mode_adj_652, tx_N_6586) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input GND_net;
    output reset_r;
    input clk_enable_28;
    input n30185;
    input n29995;
    input clk_1MHz;
    input clk_enable_178;
    input \spi_data_r[0] ;
    output n30188;
    output [39:0]spi_data_out_r_39__N_4854;
    input \spi_data_out_r_39__N_5105[0] ;
    input resetn_c;
    output \SLO_buf[0] ;
    input \spi_data_r[2] ;
    input \spi_data_r[1] ;
    output spi_data_out_r_39__N_4894;
    input spi_data_out_r_39__N_5191;
    output digital_output_r;
    input clk_enable_254;
    input n28554;
    input pin_io_c_38;
    input \spi_data_out_r_39__N_5105[1] ;
    input \spi_data_out_r_39__N_5105[2] ;
    input \spi_data_out_r_39__N_5105[3] ;
    input \spi_data_out_r_39__N_5105[4] ;
    input \spi_data_out_r_39__N_5105[5] ;
    input \spi_data_out_r_39__N_5105[6] ;
    input \spi_data_out_r_39__N_5105[7] ;
    input \spi_data_out_r_39__N_5105[8] ;
    input \spi_data_out_r_39__N_5105[9] ;
    input \spi_data_out_r_39__N_5105[10] ;
    input \spi_data_out_r_39__N_5105[11] ;
    input \spi_data_out_r_39__N_5105[12] ;
    input \spi_data_out_r_39__N_5105[13] ;
    input \spi_data_out_r_39__N_5105[14] ;
    input \spi_data_out_r_39__N_5105[15] ;
    input n29991;
    input \spi_data_out_r_39__N_5105[32] ;
    input \spi_data_out_r_39__N_5105[33] ;
    input \spi_data_out_r_39__N_5105[34] ;
    input \spi_data_out_r_39__N_5105[35] ;
    output \SLO_buf[10] ;
    output \SLO_buf[11] ;
    output \SLO_buf[12] ;
    output \SLO_buf[13] ;
    output \SLO_buf[1] ;
    output \SLO_buf[2] ;
    output \SLO_buf[3] ;
    output \SLO_buf[4] ;
    output \SLO_buf[5] ;
    output \SLO_buf[6] ;
    output \SLO_buf[7] ;
    output \SLO_buf[8] ;
    output \SLO_buf[9] ;
    output \SLO_buf[14] ;
    output \SLO_buf[15] ;
    output \SLO_buf[16] ;
    output \SLO_buf[17] ;
    output \SLO_buf[18] ;
    output \SLO_buf[19] ;
    output \SLO_buf[20] ;
    output \SLO_buf[21] ;
    output \SLO_buf[22] ;
    output \SLO_buf[23] ;
    output \SLO_buf[24] ;
    output \SLO_buf[25] ;
    output \SLO_buf[26] ;
    output \SLO_buf[27] ;
    output \SLO_buf[28] ;
    output \SLO_buf[29] ;
    output NSL;
    input \quad_homing[0] ;
    input pin_io_c_34;
    output n25873;
    input mode;
    input \cs_decoded[6] ;
    output n7170;
    output n30082;
    output n7166;
    output n30091;
    input pin_io_out_35;
    output n29943;
    input pin_io_c_33;
    output \pin_intrpt[10] ;
    input pin_io_c_32;
    output \pin_intrpt[9] ;
    output \pin_intrpt[11] ;
    output n7269;
    input UC_TXD0_c;
    output OW_ID_N_5147;
    input n30050;
    output ENC_O_N_5155;
    output OW_ID_N_5153;
    output \quad_a[3] ;
    input pin_io_out_39;
    output \quad_b[3] ;
    input \uart_slot_en[1] ;
    input \uart_slot_en[0] ;
    input n10696;
    input mode_adj_652;
    output tx_N_6586;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire clk_1MHz /* synthesis SET_AS_NETWORK=clk_1MHz, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(136[6:14])
    wire \pin_intrpt[11]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[11] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    wire [51:0]SLO;   // c:/s_links/sources/slot_cards/stepper.v(63[12:15])
    
    wire clk_enable_1134, n12344;
    wire [7:0]Cnt;   // c:/s_links/sources/slot_cards/stepper.v(62[11:14])
    
    wire clk_1MHz_enable_27;
    wire [7:0]n199;
    wire [2:0]n1;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    wire prev_MA_Temp, MA_Temp, prev_MA;
    wire [11:0]n93;
    wire [11:0]n53;
    
    wire SLO_buf_51__N_5044, clk_1MHz_enable_13, MA_Temp_N_5173, n21980;
    wire [11:0]Cnt_NSL;   // c:/s_links/sources/slot_cards/stepper.v(61[12:19])
    
    wire n21979, n21978, n30009, n28324, n30081, n28596, n28595, 
        n12089;
    wire [51:0]SLO_buf;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire n21977, n21976, n30089, n30008, NSL_N_5186, n21975, n30205, 
        n30206, n30189, n26337, n26339, n30187, n18027, clk_1MHz_enable_67, 
        n21948;
    wire [31:0]n153;
    
    wire n21947, n30186, n21946, n21945, n30204, n18025, n30088, 
        n27417, OW_ID_N_5148, n30208, n30126, n30032, n30201, n4;
    
    FD1P3IX SLO__i19 (.D(SLO[17]), .SP(clk_enable_1134), .CD(GND_net), 
            .CK(clk), .Q(SLO[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i19.GSR = "DISABLED";
    FD1P3IX SLO__i20 (.D(SLO[18]), .SP(clk_enable_1134), .CD(GND_net), 
            .CK(clk), .Q(SLO[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i20.GSR = "DISABLED";
    FD1P3IX SLO__i42 (.D(SLO[40]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i42.GSR = "DISABLED";
    FD1P3IX SLO__i21 (.D(SLO[19]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i21.GSR = "DISABLED";
    FD1P3IX SLO__i22 (.D(SLO[20]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i22.GSR = "DISABLED";
    FD1P3IX reset_r_491 (.D(n29995), .SP(clk_enable_28), .CD(n30185), 
            .CK(clk), .Q(reset_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam reset_r_491.GSR = "DISABLED";
    FD1P3IX SLO__i23 (.D(SLO[21]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i23.GSR = "DISABLED";
    FD1P3IX Cnt__i0 (.D(n199[0]), .SP(clk_1MHz_enable_27), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i0.GSR = "DISABLED";
    FD1P3IX SLO__i24 (.D(SLO[22]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i24.GSR = "DISABLED";
    FD1P3IX SLO__i25 (.D(SLO[23]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i25.GSR = "DISABLED";
    FD1P3IX SLO__i26 (.D(SLO[24]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i26.GSR = "DISABLED";
    FD1P3IX SLO__i27 (.D(SLO[25]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i27.GSR = "DISABLED";
    FD1P3IX mode__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_178), .CD(n30185), 
            .CK(clk), .Q(n1[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i0.GSR = "DISABLED";
    FD1S3AX prev_MA_Temp_487 (.D(MA_Temp), .CK(clk), .Q(prev_MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam prev_MA_Temp_487.GSR = "DISABLED";
    FD1S3AX prev_MA_489 (.D(n30188), .CK(clk), .Q(prev_MA)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam prev_MA_489.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i0 (.D(\spi_data_out_r_39__N_5105[0] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i0.GSR = "DISABLED";
    FD1P3IX SLO__i28 (.D(SLO[26]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i28.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1781__i0 (.D(n53[0]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781__i0.GSR = "DISABLED";
    FD1P3AX SLO_buf__i1 (.D(SLO[0]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i1.GSR = "DISABLED";
    FD1P3IX SLO__i29 (.D(SLO[27]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i29.GSR = "DISABLED";
    FD1P3IX mode__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_178), .CD(n30185), 
            .CK(clk), .Q(n1[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i2.GSR = "DISABLED";
    FD1P3IX mode__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_178), .CD(n30185), 
            .CK(clk), .Q(n1[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i1.GSR = "DISABLED";
    FD1P3IX SLO__i30 (.D(SLO[28]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i30.GSR = "DISABLED";
    FD1P3IX SLO__i31 (.D(SLO[29]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i31.GSR = "DISABLED";
    FD1S3IX i168_494 (.D(spi_data_out_r_39__N_5191), .CK(clk), .CD(n30185), 
            .Q(spi_data_out_r_39__N_4894)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam i168_494.GSR = "DISABLED";
    FD1P3IX digital_output_r_492 (.D(n28554), .SP(clk_enable_254), .CD(n30185), 
            .CK(clk), .Q(digital_output_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam digital_output_r_492.GSR = "DISABLED";
    FD1P3IX SLO__i32 (.D(SLO[30]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i32.GSR = "DISABLED";
    FD1P3IX SLO__i2 (.D(SLO[0]), .SP(clk_enable_1134), .CD(GND_net), .CK(clk), 
            .Q(SLO[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i2.GSR = "DISABLED";
    FD1P3IX SLO__i33 (.D(SLO[31]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i33.GSR = "DISABLED";
    FD1P3IX MA_Temp_483 (.D(MA_Temp_N_5173), .SP(clk_1MHz_enable_13), .CD(n30185), 
            .CK(clk_1MHz), .Q(MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam MA_Temp_483.GSR = "DISABLED";
    FD1P3IX SLO__i34 (.D(SLO[32]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i34.GSR = "DISABLED";
    FD1P3IX SLO__i35 (.D(SLO[33]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i35.GSR = "DISABLED";
    FD1P3IX SLO__i36 (.D(SLO[34]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i36.GSR = "DISABLED";
    CCU2D Cnt_NSL_1781_add_4_13 (.A0(Cnt_NSL[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21980), .S0(n53[11]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781_add_4_13.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1781_add_4_13.INIT1 = 16'h0000;
    defparam Cnt_NSL_1781_add_4_13.INJECT1_0 = "NO";
    defparam Cnt_NSL_1781_add_4_13.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1781_add_4_11 (.A0(Cnt_NSL[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Cnt_NSL[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21979), .COUT(n21980), .S0(n53[9]), .S1(n53[10]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781_add_4_11.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1781_add_4_11.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1781_add_4_11.INJECT1_0 = "NO";
    defparam Cnt_NSL_1781_add_4_11.INJECT1_1 = "NO";
    FD1P3IX SLO__i37 (.D(SLO[35]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i37.GSR = "DISABLED";
    CCU2D Cnt_NSL_1781_add_4_9 (.A0(Cnt_NSL[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Cnt_NSL[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21978), .COUT(n21979), .S0(n53[7]), .S1(n53[8]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781_add_4_9.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1781_add_4_9.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1781_add_4_9.INJECT1_0 = "NO";
    defparam Cnt_NSL_1781_add_4_9.INJECT1_1 = "NO";
    LUT4 i23907_1_lut_4_lut (.A(n30009), .B(MA_Temp), .C(n28324), .D(n30081), 
         .Z(n28596)) /* synthesis lut_function=(!(A+!(B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i23907_1_lut_4_lut.init = 16'h4414;
    FD1P3IX Cnt__i7 (.D(n199[7]), .SP(clk_1MHz_enable_27), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i7.GSR = "DISABLED";
    FD1P3IX Cnt__i6 (.D(n199[6]), .SP(clk_1MHz_enable_27), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i6.GSR = "DISABLED";
    FD1P3IX Cnt__i5 (.D(n199[5]), .SP(clk_1MHz_enable_27), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i5.GSR = "DISABLED";
    FD1P3IX Cnt__i4 (.D(n199[4]), .SP(clk_1MHz_enable_27), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i4.GSR = "DISABLED";
    FD1P3IX Cnt__i3 (.D(n199[3]), .SP(clk_1MHz_enable_27), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i3.GSR = "DISABLED";
    FD1P3IX Cnt__i2 (.D(n199[2]), .SP(clk_1MHz_enable_27), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i1 (.D(n199[1]), .SP(clk_1MHz_enable_27), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i1.GSR = "DISABLED";
    FD1P3IX SLO__i3 (.D(SLO[1]), .SP(clk_enable_1134), .CD(GND_net), .CK(clk), 
            .Q(SLO[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i3.GSR = "DISABLED";
    FD1P3IX SLO__i38 (.D(SLO[36]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i38.GSR = "DISABLED";
    FD1P3IX SLO__i39 (.D(SLO[37]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i39.GSR = "DISABLED";
    FD1P3IX SLO__i4 (.D(SLO[2]), .SP(clk_enable_1134), .CD(GND_net), .CK(clk), 
            .Q(SLO[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i4.GSR = "DISABLED";
    FD1P3IX SLO__i40 (.D(SLO[38]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i40.GSR = "DISABLED";
    FD1P3IX SLO__i41 (.D(SLO[39]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i41.GSR = "DISABLED";
    PFUMX i10337 (.BLUT(n28595), .ALUT(n28596), .C0(n12089), .Z(MA_Temp_N_5173));
    FD1P3IX SLO__i5 (.D(SLO[3]), .SP(clk_enable_1134), .CD(GND_net), .CK(clk), 
            .Q(SLO[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i5.GSR = "DISABLED";
    FD1P3IX SLO__i1 (.D(pin_io_c_38), .SP(clk_enable_1134), .CD(GND_net), 
            .CK(clk), .Q(SLO[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_5105[1] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_5105[2] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_5105[3] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_5105[4] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_5105[5] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_5105[6] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_5105[7] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_5105[8] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_5105[9] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_5105[10] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_5105[11] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_5105[12] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_5105[13] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_5105[14] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_5105[15] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i16 (.D(SLO_buf[30]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i17 (.D(SLO_buf[31]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i18 (.D(SLO_buf[32]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i19 (.D(SLO_buf[33]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i20 (.D(SLO_buf[34]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i21 (.D(SLO_buf[35]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i22 (.D(SLO_buf[36]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i23 (.D(SLO_buf[37]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i24 (.D(SLO_buf[38]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i25 (.D(SLO_buf[39]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i26 (.D(SLO_buf[40]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i27 (.D(SLO_buf[41]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i28 (.D(SLO_buf[42]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i29 (.D(SLO_buf[43]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i30 (.D(SLO_buf[44]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i31 (.D(SLO_buf[45]), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_5105[32] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i33 (.D(\spi_data_out_r_39__N_5105[33] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i33.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i34 (.D(\spi_data_out_r_39__N_5105[34] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i34.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i35 (.D(\spi_data_out_r_39__N_5105[35] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4854[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i35.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i36 (.D(\SLO_buf[10] ), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i36.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i37 (.D(\SLO_buf[11] ), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i37.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i38 (.D(\SLO_buf[12] ), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i38.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i39 (.D(\SLO_buf[13] ), .CK(clk), .CD(n29991), 
            .Q(spi_data_out_r_39__N_4854[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i39.GSR = "DISABLED";
    CCU2D Cnt_NSL_1781_add_4_7 (.A0(n93[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21977), .COUT(n21978), .S0(n53[5]), .S1(n53[6]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781_add_4_7.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1781_add_4_7.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1781_add_4_7.INJECT1_0 = "NO";
    defparam Cnt_NSL_1781_add_4_7.INJECT1_1 = "NO";
    FD1P3AX Cnt_NSL_1781__i1 (.D(n53[1]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781__i1.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1781__i2 (.D(n53[2]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781__i2.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1781__i3 (.D(n53[3]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781__i3.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1781__i4 (.D(n53[4]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781__i4.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1781__i5 (.D(n53[5]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781__i5.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1781__i6 (.D(n53[6]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781__i6.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1781__i7 (.D(n53[7]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781__i7.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1781__i8 (.D(n53[8]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781__i8.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1781__i9 (.D(n53[9]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781__i9.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1781__i10 (.D(n53[10]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781__i10.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1781__i11 (.D(n53[11]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781__i11.GSR = "DISABLED";
    FD1P3AX SLO_buf__i2 (.D(SLO[1]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i2.GSR = "DISABLED";
    FD1P3AX SLO_buf__i3 (.D(SLO[2]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i3.GSR = "DISABLED";
    FD1P3AX SLO_buf__i4 (.D(SLO[3]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i4.GSR = "DISABLED";
    FD1P3AX SLO_buf__i5 (.D(SLO[4]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i5.GSR = "DISABLED";
    FD1P3AX SLO_buf__i6 (.D(SLO[5]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i6.GSR = "DISABLED";
    FD1P3AX SLO_buf__i7 (.D(SLO[6]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i7.GSR = "DISABLED";
    FD1P3AX SLO_buf__i8 (.D(SLO[7]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i8.GSR = "DISABLED";
    FD1P3AX SLO_buf__i9 (.D(SLO[8]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i9.GSR = "DISABLED";
    FD1P3AX SLO_buf__i10 (.D(SLO[9]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i10.GSR = "DISABLED";
    FD1P3AX SLO_buf__i11 (.D(SLO[10]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i11.GSR = "DISABLED";
    FD1P3AX SLO_buf__i12 (.D(SLO[11]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i12.GSR = "DISABLED";
    FD1P3AX SLO_buf__i13 (.D(SLO[12]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i13.GSR = "DISABLED";
    FD1P3AX SLO_buf__i14 (.D(SLO[13]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i14.GSR = "DISABLED";
    FD1P3AX SLO_buf__i15 (.D(SLO[14]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i15.GSR = "DISABLED";
    FD1P3AX SLO_buf__i16 (.D(SLO[15]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i16.GSR = "DISABLED";
    FD1P3AX SLO_buf__i17 (.D(SLO[16]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i17.GSR = "DISABLED";
    FD1P3AX SLO_buf__i18 (.D(SLO[17]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i18.GSR = "DISABLED";
    FD1P3AX SLO_buf__i19 (.D(SLO[18]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i19.GSR = "DISABLED";
    FD1P3AX SLO_buf__i20 (.D(SLO[19]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i20.GSR = "DISABLED";
    FD1P3AX SLO_buf__i21 (.D(SLO[20]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i21.GSR = "DISABLED";
    FD1P3AX SLO_buf__i22 (.D(SLO[21]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i22.GSR = "DISABLED";
    FD1P3AX SLO_buf__i23 (.D(SLO[22]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i23.GSR = "DISABLED";
    FD1P3AX SLO_buf__i24 (.D(SLO[23]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i24.GSR = "DISABLED";
    FD1P3AX SLO_buf__i25 (.D(SLO[24]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i25.GSR = "DISABLED";
    FD1P3AX SLO_buf__i26 (.D(SLO[25]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i26.GSR = "DISABLED";
    FD1P3AX SLO_buf__i27 (.D(SLO[26]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i27.GSR = "DISABLED";
    FD1P3AX SLO_buf__i28 (.D(SLO[27]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i28.GSR = "DISABLED";
    FD1P3AX SLO_buf__i29 (.D(SLO[28]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i29.GSR = "DISABLED";
    FD1P3AX SLO_buf__i30 (.D(SLO[29]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(\SLO_buf[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i30.GSR = "DISABLED";
    FD1P3AX SLO_buf__i31 (.D(SLO[30]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i31.GSR = "DISABLED";
    FD1P3AX SLO_buf__i32 (.D(SLO[31]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i32.GSR = "DISABLED";
    FD1P3AX SLO_buf__i33 (.D(SLO[32]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i33.GSR = "DISABLED";
    FD1P3AX SLO_buf__i34 (.D(SLO[33]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i34.GSR = "DISABLED";
    FD1P3AX SLO_buf__i35 (.D(SLO[34]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i35.GSR = "DISABLED";
    FD1P3AX SLO_buf__i36 (.D(SLO[35]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i36.GSR = "DISABLED";
    FD1P3AX SLO_buf__i37 (.D(SLO[36]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i37.GSR = "DISABLED";
    FD1P3AX SLO_buf__i38 (.D(SLO[37]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i38.GSR = "DISABLED";
    FD1P3AX SLO_buf__i39 (.D(SLO[38]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i39.GSR = "DISABLED";
    FD1P3AX SLO_buf__i40 (.D(SLO[39]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i40.GSR = "DISABLED";
    FD1P3AX SLO_buf__i41 (.D(SLO[40]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i41.GSR = "DISABLED";
    FD1P3AX SLO_buf__i42 (.D(SLO[41]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i42.GSR = "DISABLED";
    FD1P3AX SLO_buf__i43 (.D(SLO[42]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i43.GSR = "DISABLED";
    FD1P3AX SLO_buf__i44 (.D(SLO[43]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i44.GSR = "DISABLED";
    FD1P3AX SLO_buf__i45 (.D(SLO[44]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i45.GSR = "DISABLED";
    FD1P3AX SLO_buf__i46 (.D(SLO[45]), .SP(SLO_buf_51__N_5044), .CK(clk), 
            .Q(SLO_buf[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i46.GSR = "DISABLED";
    FD1P3IX SLO__i6 (.D(SLO[4]), .SP(clk_enable_1134), .CD(GND_net), .CK(clk), 
            .Q(SLO[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i6.GSR = "DISABLED";
    CCU2D Cnt_NSL_1781_add_4_5 (.A0(n93[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21976), .COUT(n21977), .S0(n53[3]), .S1(n53[4]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781_add_4_5.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1781_add_4_5.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1781_add_4_5.INJECT1_0 = "NO";
    defparam Cnt_NSL_1781_add_4_5.INJECT1_1 = "NO";
    LUT4 SLO_buf_51__I_166_2_lut (.A(prev_MA_Temp), .B(MA_Temp), .Z(SLO_buf_51__N_5044)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[5:38])
    defparam SLO_buf_51__I_166_2_lut.init = 16'h2222;
    LUT4 i23975_4_lut (.A(NSL), .B(n30089), .C(n12089), .D(n30008), 
         .Z(NSL_N_5186)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C+(D))))) */ ;
    defparam i23975_4_lut.init = 16'h3b37;
    CCU2D Cnt_NSL_1781_add_4_3 (.A0(n93[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21975), .COUT(n21976), .S0(n53[1]), .S1(n53[2]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781_add_4_3.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1781_add_4_3.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1781_add_4_3.INJECT1_0 = "NO";
    defparam Cnt_NSL_1781_add_4_3.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1781_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n30205), .B1(n30206), .C1(n93[0]), .D1(GND_net), 
          .COUT(n21975), .S1(n53[0]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1781_add_4_1.INIT0 = 16'hF000;
    defparam Cnt_NSL_1781_add_4_1.INIT1 = 16'h8787;
    defparam Cnt_NSL_1781_add_4_1.INJECT1_0 = "NO";
    defparam Cnt_NSL_1781_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(\quad_homing[0] ), .B(pin_io_c_34), .Z(n25873)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(74[8:17])
    defparam i1_2_lut.init = 16'h8888;
    FD1P3IX SLO__i7 (.D(SLO[5]), .SP(clk_enable_1134), .CD(GND_net), .CK(clk), 
            .Q(SLO[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i7.GSR = "DISABLED";
    LUT4 i24153_4_lut_4_lut (.A(n1[2]), .B(n30189), .C(n26337), .D(n26339), 
         .Z(clk_enable_1134)) /* synthesis lut_function=(!(A (B+(D))+!A ((D)+!C))) */ ;
    defparam i24153_4_lut_4_lut.init = 16'h0072;
    LUT4 Select_2832_i3_3_lut_4_lut (.A(n1[2]), .B(n30189), .C(mode), 
         .D(\cs_decoded[6] ), .Z(n7170)) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;
    defparam Select_2832_i3_3_lut_4_lut.init = 16'hf222;
    LUT4 i13705_2_lut_4_lut (.A(Cnt[1]), .B(n30187), .C(Cnt[0]), .D(Cnt[4]), 
         .Z(n18027)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam i13705_2_lut_4_lut.init = 16'hec00;
    LUT4 i24162_3_lut_4_lut (.A(n30206), .B(n30205), .C(n12089), .D(resetn_c), 
         .Z(clk_1MHz_enable_67)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i24162_3_lut_4_lut.init = 16'h7f00;
    CCU2D add_564_9 (.A0(Cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21948), 
          .S0(n153[7]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_9.INIT0 = 16'h5aaa;
    defparam add_564_9.INIT1 = 16'h0000;
    defparam add_564_9.INJECT1_0 = "NO";
    defparam add_564_9.INJECT1_1 = "NO";
    CCU2D add_564_7 (.A0(Cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21947), 
          .COUT(n21948), .S0(n153[5]), .S1(n153[6]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_7.INIT0 = 16'h5aaa;
    defparam add_564_7.INIT1 = 16'h5aaa;
    defparam add_564_7.INJECT1_0 = "NO";
    defparam add_564_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(n30186), .B(n18027), .C(Cnt[5]), .D(n30082), .Z(n12089)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut.init = 16'hfffe;
    CCU2D add_564_5 (.A0(Cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21946), 
          .COUT(n21947), .S0(n153[3]), .S1(n153[4]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_5.INIT0 = 16'h5aaa;
    defparam add_564_5.INIT1 = 16'h5aaa;
    defparam add_564_5.INJECT1_0 = "NO";
    defparam add_564_5.INJECT1_1 = "NO";
    CCU2D add_564_3 (.A0(Cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21945), 
          .COUT(n21946), .S0(n153[1]), .S1(n153[2]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_3.INIT0 = 16'h5aaa;
    defparam add_564_3.INIT1 = 16'h5aaa;
    defparam add_564_3.INJECT1_0 = "NO";
    defparam add_564_3.INJECT1_1 = "NO";
    CCU2D add_564_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n21945), 
          .S1(n153[0]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_1.INIT0 = 16'hF000;
    defparam add_564_1.INIT1 = 16'h5555;
    defparam add_564_1.INJECT1_0 = "NO";
    defparam add_564_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_786 (.A(Cnt[6]), .B(Cnt[7]), .Z(n30186)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_786.init = 16'heeee;
    LUT4 i1_3_lut_rep_681_4_lut (.A(Cnt[6]), .B(Cnt[7]), .C(Cnt[0]), .D(n30187), 
         .Z(n30081)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_rep_681_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut (.A(Cnt[6]), .B(Cnt[7]), .C(n1[0]), .D(n30204), 
         .Z(n18025)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hffef;
    LUT4 i1_2_lut_rep_787 (.A(Cnt[2]), .B(Cnt[3]), .Z(n30187)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_787.init = 16'heeee;
    LUT4 i1_3_lut_rep_688_4_lut (.A(Cnt[2]), .B(Cnt[3]), .C(Cnt[0]), .D(Cnt[1]), 
         .Z(n30088)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_3_lut_rep_688_4_lut.init = 16'hfeee;
    LUT4 i23979_2_lut_rep_788 (.A(MA_Temp), .B(clk_1MHz), .Z(n30188)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i23979_2_lut_rep_788.init = 16'h7777;
    LUT4 i1_2_lut_3_lut (.A(MA_Temp), .B(clk_1MHz), .C(prev_MA), .Z(n26339)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_3_lut_adj_820 (.A(MA_Temp), .B(clk_1MHz), .C(n1[2]), 
         .Z(n27417)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i1_2_lut_3_lut_adj_820.init = 16'h7070;
    LUT4 i1_2_lut_rep_789 (.A(n1[0]), .B(n1[1]), .Z(n30189)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_789.init = 16'heeee;
    LUT4 i1_2_lut_rep_682_3_lut (.A(n1[0]), .B(n1[1]), .C(n1[2]), .Z(n30082)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_rep_682_3_lut.init = 16'hefef;
    LUT4 i24037_2_lut_3_lut_4_lut (.A(n1[0]), .B(n1[1]), .C(mode), .D(n1[2]), 
         .Z(n7166)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+(D))))) */ ;
    defparam i24037_2_lut_3_lut_4_lut.init = 16'h0e0f;
    LUT4 i1_2_lut_rep_691_3_lut (.A(n1[0]), .B(n1[1]), .C(n1[2]), .Z(n30091)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_691_3_lut.init = 16'hfefe;
    LUT4 RESET_N_4460_bdd_2_lut_24382_3_lut_4_lut (.A(n1[0]), .B(n1[1]), 
         .C(pin_io_out_35), .D(n1[2]), .Z(n29943)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam RESET_N_4460_bdd_2_lut_24382_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2980_2_lut_3_lut_4_lut (.A(n1[0]), .B(n1[1]), .C(pin_io_c_33), 
         .D(n1[2]), .Z(\pin_intrpt[10] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i2980_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2979_2_lut_3_lut_4_lut (.A(n1[0]), .B(n1[1]), .C(pin_io_c_32), 
         .D(n1[2]), .Z(\pin_intrpt[9] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i2979_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2981_2_lut_3_lut_4_lut (.A(n1[0]), .B(n1[1]), .C(pin_io_c_34), 
         .D(n1[2]), .Z(\pin_intrpt[11] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i2981_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2955_1_lut_2_lut_3_lut (.A(n1[0]), .B(n1[1]), .C(n1[2]), .Z(n7269)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i2955_1_lut_2_lut_3_lut.init = 16'h0101;
    LUT4 digital_output_r_I_0_547_3_lut (.A(digital_output_r), .B(UC_TXD0_c), 
         .C(OW_ID_N_5148), .Z(OW_ID_N_5147)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[16] 91[59])
    defparam digital_output_r_I_0_547_3_lut.init = 16'hcaca;
    LUT4 i4_4_lut (.A(n30208), .B(n30050), .C(n30126), .D(n1[0]), .Z(OW_ID_N_5148)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i4_4_lut.init = 16'h4000;
    LUT4 i24079_3_lut (.A(n1[0]), .B(n1[2]), .C(n1[1]), .Z(ENC_O_N_5155)) /* synthesis lut_function=(!(A (B+(C))+!A (B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(80[8:13])
    defparam i24079_3_lut.init = 16'h1313;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n30032), .B(n18025), .C(n153[0]), .D(n12089), 
         .Z(n199[0])) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h10f0;
    LUT4 i13673_2_lut_rep_801 (.A(Cnt[1]), .B(Cnt[4]), .Z(n30201)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13673_2_lut_rep_801.init = 16'h8888;
    LUT4 i23622_2_lut_3_lut (.A(Cnt[1]), .B(Cnt[4]), .C(Cnt[5]), .Z(n28324)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i23622_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_608_3_lut_4_lut (.A(Cnt[1]), .B(Cnt[4]), .C(n30081), 
         .D(Cnt[5]), .Z(n30008)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_rep_608_3_lut_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut_3_lut_4_lut_adj_821 (.A(n30032), .B(n18025), .C(n153[7]), 
         .D(n12089), .Z(n199[7])) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_821.init = 16'h10f0;
    LUT4 i1_2_lut_rep_804 (.A(n1[2]), .B(n1[1]), .Z(n30204)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i1_2_lut_rep_804.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_4_lut_adj_822 (.A(n30032), .B(n18025), .C(n153[6]), 
         .D(n12089), .Z(n199[6])) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_822.init = 16'h10f0;
    LUT4 i24076_3_lut_4_lut (.A(n1[2]), .B(n1[1]), .C(n1[0]), .D(OW_ID_N_5148), 
         .Z(OW_ID_N_5153)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i24076_3_lut_4_lut.init = 16'h00fb;
    LUT4 i1_3_lut_rep_805 (.A(Cnt_NSL[9]), .B(Cnt_NSL[8]), .C(Cnt_NSL[7]), 
         .Z(n30205)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_rep_805.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut_adj_823 (.A(n30032), .B(n18025), .C(n153[5]), 
         .D(n12089), .Z(n199[5])) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_823.init = 16'h10f0;
    LUT4 i1_2_lut_rep_689_4_lut (.A(Cnt_NSL[9]), .B(Cnt_NSL[8]), .C(Cnt_NSL[7]), 
         .D(n30206), .Z(n30089)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_rep_689_4_lut.init = 16'hfe00;
    LUT4 i1_2_lut_rep_806 (.A(Cnt_NSL[11]), .B(Cnt_NSL[10]), .Z(n30206)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i1_2_lut_rep_806.init = 16'h8888;
    LUT4 i24165_2_lut_3_lut_4_lut (.A(Cnt_NSL[11]), .B(Cnt_NSL[10]), .C(resetn_c), 
         .D(n30205), .Z(clk_1MHz_enable_27)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i24165_2_lut_3_lut_4_lut.init = 16'h8f0f;
    LUT4 i1_2_lut_3_lut_4_lut_adj_824 (.A(n30032), .B(n18025), .C(n153[4]), 
         .D(n12089), .Z(n199[4])) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_824.init = 16'h10f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_825 (.A(n30032), .B(n18025), .C(n153[3]), 
         .D(n12089), .Z(n199[3])) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_825.init = 16'h10f0;
    LUT4 i1_2_lut_rep_808 (.A(n1[2]), .B(n1[1]), .Z(n30208)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i1_2_lut_rep_808.init = 16'heeee;
    LUT4 i2982_2_lut_3_lut_4_lut (.A(n1[2]), .B(n1[1]), .C(pin_io_c_38), 
         .D(n1[0]), .Z(\quad_a[3] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i2982_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i2983_2_lut_3_lut_4_lut (.A(n1[2]), .B(n1[1]), .C(pin_io_out_39), 
         .D(n1[0]), .Z(\quad_b[3] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i2983_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_826 (.A(n30032), .B(n18025), .C(n153[2]), 
         .D(n12089), .Z(n199[2])) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_826.init = 16'h10f0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_827 (.A(n30032), .B(n18025), .C(n153[1]), 
         .D(n12089), .Z(n199[1])) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_827.init = 16'h10f0;
    LUT4 i24167_4_lut (.A(clk_1MHz_enable_27), .B(n30032), .C(n12089), 
         .D(n18025), .Z(clk_1MHz_enable_13)) /* synthesis lut_function=(!((B (C+!(D))+!B (C (D)))+!A)) */ ;
    defparam i24167_4_lut.init = 16'h0a22;
    LUT4 i1_4_lut_adj_828 (.A(n1[1]), .B(n1[0]), .C(Cnt[1]), .D(n4), 
         .Z(n26337)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_828.init = 16'h8880;
    LUT4 i1_2_lut_3_lut_adj_829 (.A(Cnt[5]), .B(n30081), .C(Cnt[4]), .Z(n4)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(133[16:19])
    defparam i1_2_lut_3_lut_adj_829.init = 16'hfefe;
    LUT4 i23906_1_lut_2_lut_3_lut_4_lut (.A(Cnt[5]), .B(n30081), .C(MA_Temp), 
         .D(n30201), .Z(n28595)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(133[16:19])
    defparam i23906_1_lut_2_lut_3_lut_4_lut.init = 16'he1f0;
    LUT4 i1_3_lut_rep_632 (.A(Cnt[4]), .B(n30088), .C(Cnt[5]), .Z(n30032)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam i1_3_lut_rep_632.init = 16'h8080;
    LUT4 i13711_2_lut_rep_609_4_lut (.A(Cnt[4]), .B(n30088), .C(Cnt[5]), 
         .D(n18025), .Z(n30009)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam i13711_2_lut_rep_609_4_lut.init = 16'hff80;
    LUT4 i1_4_lut_adj_830 (.A(n1[0]), .B(n1[1]), .C(prev_MA), .D(n27417), 
         .Z(n12344)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_830.init = 16'h0100;
    FD1P3AX NSL_484 (.D(NSL_N_5186), .SP(clk_1MHz_enable_67), .CK(clk_1MHz), 
            .Q(NSL)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam NSL_484.GSR = "DISABLED";
    FD1P3IX SLO__i8 (.D(SLO[6]), .SP(clk_enable_1134), .CD(GND_net), .CK(clk), 
            .Q(SLO[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i8.GSR = "DISABLED";
    FD1P3IX SLO__i9 (.D(SLO[7]), .SP(clk_enable_1134), .CD(GND_net), .CK(clk), 
            .Q(SLO[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i9.GSR = "DISABLED";
    FD1P3IX SLO__i10 (.D(SLO[8]), .SP(clk_enable_1134), .CD(GND_net), 
            .CK(clk), .Q(SLO[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i10.GSR = "DISABLED";
    FD1P3IX SLO__i11 (.D(SLO[9]), .SP(clk_enable_1134), .CD(GND_net), 
            .CK(clk), .Q(SLO[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i11.GSR = "DISABLED";
    FD1P3IX SLO__i43 (.D(SLO[41]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i43.GSR = "DISABLED";
    FD1P3IX SLO__i44 (.D(SLO[42]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i44.GSR = "DISABLED";
    FD1P3IX SLO__i12 (.D(SLO[10]), .SP(clk_enable_1134), .CD(GND_net), 
            .CK(clk), .Q(SLO[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i12.GSR = "DISABLED";
    FD1P3IX SLO__i13 (.D(SLO[11]), .SP(clk_enable_1134), .CD(GND_net), 
            .CK(clk), .Q(SLO[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i13.GSR = "DISABLED";
    FD1P3IX SLO__i14 (.D(SLO[12]), .SP(clk_enable_1134), .CD(GND_net), 
            .CK(clk), .Q(SLO[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i14.GSR = "DISABLED";
    FD1P3IX SLO__i46 (.D(SLO[44]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i46.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_726 (.A(\uart_slot_en[1] ), .B(\uart_slot_en[0] ), 
         .Z(n30126)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_726.init = 16'h2222;
    FD1P3IX SLO__i45 (.D(SLO[43]), .SP(clk_enable_1134), .CD(n12344), 
            .CK(clk), .Q(SLO[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i45.GSR = "DISABLED";
    LUT4 i24032_3_lut_4_lut (.A(\uart_slot_en[1] ), .B(\uart_slot_en[0] ), 
         .C(n10696), .D(mode_adj_652), .Z(tx_N_6586)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;
    defparam i24032_3_lut_4_lut.init = 16'hdfff;
    FD1P3IX SLO__i15 (.D(SLO[13]), .SP(clk_enable_1134), .CD(GND_net), 
            .CK(clk), .Q(SLO[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i15.GSR = "DISABLED";
    FD1P3IX SLO__i16 (.D(SLO[14]), .SP(clk_enable_1134), .CD(GND_net), 
            .CK(clk), .Q(SLO[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i16.GSR = "DISABLED";
    FD1P3IX SLO__i17 (.D(SLO[15]), .SP(clk_enable_1134), .CD(GND_net), 
            .CK(clk), .Q(SLO[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i17.GSR = "DISABLED";
    FD1P3IX SLO__i18 (.D(SLO[16]), .SP(clk_enable_1134), .CD(GND_net), 
            .CK(clk), .Q(SLO[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i18.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \stepper(DEV_ID=4,UART_ADDRESS_WIDTH=4) 
//

module \stepper(DEV_ID=4,UART_ADDRESS_WIDTH=4)  (reset_r, clk, n30185, 
            n30031, clk_1MHz, GND_net, n30146, clk_enable_641, \spi_data_r[0] , 
            spi_data_out_r_39__N_5197, resetn_c, digital_output_r, n28549, 
            \uart_slot_en[0] , n30091, n29594, spi_data_out_r_39__N_5237, 
            spi_data_out_r_39__N_5534, pin_io_out_45, \uart_slot_en[2] , 
            n29481, pin_io_c_48, \spi_data_r[1] , \spi_data_r[2] , n47, 
            NSL, n25979, n23916, n30199, \quad_homing[0] , pin_io_c_44, 
            n25893, ENC_O_N_5498, n30180, TX_IN_N_6565, n7163, \uart_slot_en[1] , 
            n23722, EM_STOP, n25699, UC_TXD0_c, OW_ID_N_5490, n30050, 
            n30120, pin_io_out_49, \quad_b[4] , \quad_a[4] , \pin_intrpt[14] , 
            n30055, OW_ID_N_5496, n7266, pin_io_c_42, \pin_intrpt[12] , 
            pin_io_c_43, \pin_intrpt[13] ) /* synthesis syn_module_defined=1 */ ;
    output reset_r;
    input clk;
    input n30185;
    input n30031;
    input clk_1MHz;
    input GND_net;
    output n30146;
    input clk_enable_641;
    input \spi_data_r[0] ;
    output [39:0]spi_data_out_r_39__N_5197;
    input resetn_c;
    output digital_output_r;
    input n28549;
    input \uart_slot_en[0] ;
    input n30091;
    output n29594;
    output spi_data_out_r_39__N_5237;
    input spi_data_out_r_39__N_5534;
    input pin_io_out_45;
    input \uart_slot_en[2] ;
    output n29481;
    input pin_io_c_48;
    input \spi_data_r[1] ;
    input \spi_data_r[2] ;
    input n47;
    output NSL;
    input n25979;
    input n23916;
    input n30199;
    input \quad_homing[0] ;
    input pin_io_c_44;
    output n25893;
    output ENC_O_N_5498;
    output n30180;
    input TX_IN_N_6565;
    output n7163;
    input \uart_slot_en[1] ;
    output n23722;
    input EM_STOP;
    input n25699;
    input UC_TXD0_c;
    output OW_ID_N_5490;
    input n30050;
    input n30120;
    input pin_io_out_49;
    output \quad_b[4] ;
    output \quad_a[4] ;
    output \pin_intrpt[14] ;
    output n30055;
    output OW_ID_N_5496;
    output n7266;
    input pin_io_c_42;
    output \pin_intrpt[12] ;
    input pin_io_c_43;
    output \pin_intrpt[13] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire clk_1MHz /* synthesis SET_AS_NETWORK=clk_1MHz, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(136[6:14])
    wire \pin_intrpt[14]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[14] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    
    wire clk_enable_36;
    wire [51:0]SLO_buf;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire SLO_buf_51__N_5387;
    wire [51:0]SLO;   // c:/s_links/sources/slot_cards/stepper.v(63[12:15])
    wire [7:0]Cnt;   // c:/s_links/sources/slot_cards/stepper.v(62[11:14])
    
    wire clk_1MHz_enable_20;
    wire [7:0]n199;
    
    wire MA_Temp, clk_1MHz_enable_8, MA_Temp_N_5516, n21993;
    wire [11:0]Cnt_NSL;   // c:/s_links/sources/slot_cards/stepper.v(61[12:19])
    wire [11:0]n53;
    
    wire prev_MA_Temp, n21992, n21991, n21990;
    wire [11:0]n93;
    
    wire n23598, n24570, n30179;
    wire [2:0]mode;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    wire n18530, n18498, n26301, n18592, prev_MA;
    wire [39:0]spi_data_out_r_39__N_5448;
    
    wire n21989, clk_enable_221, n21988, n30128, n30183, n30184, 
        clk_enable_1103, n28589, n28590, n30079, n30002, NSL_N_5529, 
        clk_1MHz_enable_68, n21959;
    wire [31:0]n153;
    
    wire n21958, n21957, n21956, n30085, n30086, n26387, n4, OW_ID_N_5491, 
        n30207, n30148, n28322, n12496;
    
    FD1P3IX reset_r_491 (.D(n30031), .SP(clk_enable_36), .CD(n30185), 
            .CK(clk), .Q(reset_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam reset_r_491.GSR = "DISABLED";
    FD1P3AX SLO_buf__i1 (.D(SLO[0]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i1.GSR = "DISABLED";
    FD1P3IX Cnt__i0 (.D(n199[0]), .SP(clk_1MHz_enable_20), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i0.GSR = "DISABLED";
    FD1P3IX MA_Temp_483 (.D(MA_Temp_N_5516), .SP(clk_1MHz_enable_8), .CD(n30185), 
            .CK(clk_1MHz), .Q(MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam MA_Temp_483.GSR = "DISABLED";
    CCU2D Cnt_NSL_1782_add_4_13 (.A0(Cnt_NSL[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21993), .S0(n53[11]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782_add_4_13.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1782_add_4_13.INIT1 = 16'h0000;
    defparam Cnt_NSL_1782_add_4_13.INJECT1_0 = "NO";
    defparam Cnt_NSL_1782_add_4_13.INJECT1_1 = "NO";
    LUT4 SLO_buf_51__I_190_2_lut (.A(prev_MA_Temp), .B(MA_Temp), .Z(SLO_buf_51__N_5387)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[5:38])
    defparam SLO_buf_51__I_190_2_lut.init = 16'h2222;
    CCU2D Cnt_NSL_1782_add_4_11 (.A0(Cnt_NSL[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Cnt_NSL[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21992), .COUT(n21993), .S0(n53[9]), .S1(n53[10]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782_add_4_11.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1782_add_4_11.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1782_add_4_11.INJECT1_0 = "NO";
    defparam Cnt_NSL_1782_add_4_11.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1782_add_4_9 (.A0(Cnt_NSL[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Cnt_NSL[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21991), .COUT(n21992), .S0(n53[7]), .S1(n53[8]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782_add_4_9.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1782_add_4_9.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1782_add_4_9.INJECT1_0 = "NO";
    defparam Cnt_NSL_1782_add_4_9.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1782_add_4_7 (.A0(n93[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21990), .COUT(n21991), .S0(n53[5]), .S1(n53[6]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782_add_4_7.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1782_add_4_7.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1782_add_4_7.INJECT1_0 = "NO";
    defparam Cnt_NSL_1782_add_4_7.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(n23598), .B(n24570), .C(n30179), .D(mode[2]), 
         .Z(n18530)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i1_4_lut.init = 16'hffef;
    FD1S3AX prev_MA_Temp_487 (.D(MA_Temp), .CK(clk), .Q(prev_MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam prev_MA_Temp_487.GSR = "DISABLED";
    LUT4 i1_3_lut (.A(Cnt[5]), .B(n18498), .C(Cnt[4]), .Z(n24570)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_adj_816 (.A(n23598), .B(n18498), .C(n26301), .D(Cnt[4]), 
         .Z(n18592)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_816.init = 16'hfefa;
    FD1S3AX prev_MA_489 (.D(n30146), .CK(clk), .Q(prev_MA)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam prev_MA_489.GSR = "DISABLED";
    FD1P3IX mode__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_641), .CD(n30185), 
            .CK(clk), .Q(mode[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i0 (.D(spi_data_out_r_39__N_5448[0]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i0.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(Cnt[6]), .B(Cnt[7]), .Z(n23598)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(109[8:17])
    defparam i1_2_lut.init = 16'heeee;
    FD1P3AX Cnt_NSL_1782__i0 (.D(n53[0]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782__i0.GSR = "DISABLED";
    CCU2D Cnt_NSL_1782_add_4_5 (.A0(n93[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21989), .COUT(n21990), .S0(n53[3]), .S1(n53[4]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782_add_4_5.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1782_add_4_5.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1782_add_4_5.INJECT1_0 = "NO";
    defparam Cnt_NSL_1782_add_4_5.INJECT1_1 = "NO";
    FD1P3IX digital_output_r_492 (.D(n28549), .SP(clk_enable_221), .CD(n30185), 
            .CK(clk), .Q(digital_output_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam digital_output_r_492.GSR = "DISABLED";
    CCU2D Cnt_NSL_1782_add_4_3 (.A0(n93[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21988), .COUT(n21989), .S0(n53[1]), .S1(n53[2]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782_add_4_3.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1782_add_4_3.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1782_add_4_3.INJECT1_0 = "NO";
    defparam Cnt_NSL_1782_add_4_3.INJECT1_1 = "NO";
    LUT4 n28_bdd_3_lut_24359_4_lut (.A(mode[1]), .B(n30128), .C(\uart_slot_en[0] ), 
         .D(n30091), .Z(n29594)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam n28_bdd_3_lut_24359_4_lut.init = 16'hefe0;
    FD1S3IX i168_494 (.D(spi_data_out_r_39__N_5534), .CK(clk), .CD(n30185), 
            .Q(spi_data_out_r_39__N_5237)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam i168_494.GSR = "DISABLED";
    LUT4 RESET_N_5489_bdd_3_lut_4_lut (.A(mode[1]), .B(n30128), .C(pin_io_out_45), 
         .D(\uart_slot_en[2] ), .Z(n29481)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam RESET_N_5489_bdd_3_lut_4_lut.init = 16'h00e0;
    CCU2D Cnt_NSL_1782_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n30183), .B1(n30184), .C1(n93[0]), .D1(GND_net), 
          .COUT(n21988), .S1(n53[0]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782_add_4_1.INIT0 = 16'hF000;
    defparam Cnt_NSL_1782_add_4_1.INIT1 = 16'h8787;
    defparam Cnt_NSL_1782_add_4_1.INJECT1_0 = "NO";
    defparam Cnt_NSL_1782_add_4_1.INJECT1_1 = "NO";
    FD1P3IX Cnt__i7 (.D(n199[7]), .SP(clk_1MHz_enable_20), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i7.GSR = "DISABLED";
    FD1P3IX Cnt__i6 (.D(n199[6]), .SP(clk_1MHz_enable_20), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i6.GSR = "DISABLED";
    FD1P3IX Cnt__i5 (.D(n199[5]), .SP(clk_1MHz_enable_20), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i5.GSR = "DISABLED";
    FD1P3IX Cnt__i4 (.D(n199[4]), .SP(clk_1MHz_enable_20), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i4.GSR = "DISABLED";
    FD1P3IX Cnt__i3 (.D(n199[3]), .SP(clk_1MHz_enable_20), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i3.GSR = "DISABLED";
    FD1P3IX Cnt__i2 (.D(n199[2]), .SP(clk_1MHz_enable_20), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i1 (.D(n199[1]), .SP(clk_1MHz_enable_20), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i1.GSR = "DISABLED";
    FD1P3AX SLO_buf__i46 (.D(SLO[45]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i46.GSR = "DISABLED";
    FD1P3AX SLO_buf__i45 (.D(SLO[44]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i45.GSR = "DISABLED";
    FD1P3AX SLO_buf__i44 (.D(SLO[43]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i44.GSR = "DISABLED";
    FD1P3AX SLO_buf__i43 (.D(SLO[42]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i43.GSR = "DISABLED";
    FD1P3AX SLO_buf__i42 (.D(SLO[41]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i42.GSR = "DISABLED";
    FD1P3AX SLO_buf__i41 (.D(SLO[40]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i41.GSR = "DISABLED";
    FD1P3AX SLO_buf__i40 (.D(SLO[39]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i40.GSR = "DISABLED";
    FD1P3AX SLO_buf__i39 (.D(SLO[38]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i39.GSR = "DISABLED";
    FD1P3AX SLO_buf__i38 (.D(SLO[37]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i38.GSR = "DISABLED";
    FD1P3AX SLO_buf__i37 (.D(SLO[36]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i37.GSR = "DISABLED";
    FD1P3AX SLO_buf__i36 (.D(SLO[35]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i36.GSR = "DISABLED";
    FD1P3AX SLO_buf__i35 (.D(SLO[34]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i35.GSR = "DISABLED";
    FD1P3AX SLO_buf__i34 (.D(SLO[33]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i34.GSR = "DISABLED";
    FD1P3AX SLO_buf__i33 (.D(SLO[32]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i33.GSR = "DISABLED";
    FD1P3AX SLO_buf__i32 (.D(SLO[31]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i32.GSR = "DISABLED";
    FD1P3AX SLO_buf__i31 (.D(SLO[30]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i31.GSR = "DISABLED";
    FD1P3AX SLO_buf__i30 (.D(SLO[29]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i30.GSR = "DISABLED";
    FD1P3AX SLO_buf__i29 (.D(SLO[28]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i29.GSR = "DISABLED";
    FD1P3AX SLO_buf__i28 (.D(SLO[27]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i28.GSR = "DISABLED";
    FD1P3AX SLO_buf__i27 (.D(SLO[26]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i27.GSR = "DISABLED";
    FD1P3AX SLO_buf__i26 (.D(SLO[25]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i26.GSR = "DISABLED";
    FD1P3AX SLO_buf__i25 (.D(SLO[24]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i25.GSR = "DISABLED";
    FD1P3AX SLO_buf__i24 (.D(SLO[23]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i24.GSR = "DISABLED";
    FD1P3AX SLO_buf__i23 (.D(SLO[22]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i23.GSR = "DISABLED";
    FD1P3AX SLO_buf__i22 (.D(SLO[21]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i22.GSR = "DISABLED";
    FD1P3AX SLO_buf__i21 (.D(SLO[20]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i21.GSR = "DISABLED";
    FD1P3AX SLO_buf__i20 (.D(SLO[19]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i20.GSR = "DISABLED";
    FD1P3AX SLO_buf__i19 (.D(SLO[18]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i19.GSR = "DISABLED";
    FD1P3AX SLO_buf__i18 (.D(SLO[17]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i18.GSR = "DISABLED";
    FD1P3AX SLO_buf__i17 (.D(SLO[16]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i17.GSR = "DISABLED";
    FD1P3AX SLO_buf__i16 (.D(SLO[15]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i16.GSR = "DISABLED";
    FD1P3AX SLO_buf__i15 (.D(SLO[14]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i15.GSR = "DISABLED";
    FD1P3AX SLO_buf__i14 (.D(SLO[13]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i14.GSR = "DISABLED";
    FD1P3AX SLO_buf__i13 (.D(SLO[12]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i13.GSR = "DISABLED";
    FD1P3AX SLO_buf__i12 (.D(SLO[11]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i12.GSR = "DISABLED";
    FD1P3AX SLO_buf__i11 (.D(SLO[10]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i11.GSR = "DISABLED";
    FD1P3AX SLO_buf__i10 (.D(SLO[9]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i10.GSR = "DISABLED";
    FD1P3AX SLO_buf__i9 (.D(SLO[8]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i9.GSR = "DISABLED";
    FD1P3AX SLO_buf__i8 (.D(SLO[7]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i8.GSR = "DISABLED";
    FD1P3AX SLO_buf__i7 (.D(SLO[6]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i7.GSR = "DISABLED";
    FD1P3AX SLO_buf__i6 (.D(SLO[5]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i6.GSR = "DISABLED";
    FD1P3AX SLO_buf__i5 (.D(SLO[4]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i5.GSR = "DISABLED";
    FD1P3AX SLO_buf__i4 (.D(SLO[3]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i4.GSR = "DISABLED";
    FD1P3AX SLO_buf__i3 (.D(SLO[2]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i3.GSR = "DISABLED";
    FD1P3AX SLO_buf__i2 (.D(SLO[1]), .SP(SLO_buf_51__N_5387), .CK(clk), 
            .Q(SLO_buf[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i2.GSR = "DISABLED";
    FD1P3IX SLO__i1 (.D(pin_io_c_48), .SP(clk_enable_1103), .CD(GND_net), 
            .CK(clk), .Q(SLO[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i1.GSR = "DISABLED";
    FD1P3IX mode__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_641), .CD(n30185), 
            .CK(clk), .Q(mode[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i1.GSR = "DISABLED";
    FD1P3IX mode__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_641), .CD(n30185), 
            .CK(clk), .Q(mode[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i2.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(spi_data_out_r_39__N_5448[1]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(spi_data_out_r_39__N_5448[2]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(spi_data_out_r_39__N_5448[3]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(spi_data_out_r_39__N_5448[4]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(spi_data_out_r_39__N_5448[5]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(spi_data_out_r_39__N_5448[6]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(spi_data_out_r_39__N_5448[7]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(spi_data_out_r_39__N_5448[8]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(spi_data_out_r_39__N_5448[9]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(spi_data_out_r_39__N_5448[10]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(spi_data_out_r_39__N_5448[11]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(spi_data_out_r_39__N_5448[12]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(spi_data_out_r_39__N_5448[13]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(spi_data_out_r_39__N_5448[14]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(spi_data_out_r_39__N_5448[15]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i16 (.D(SLO_buf[30]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i17 (.D(SLO_buf[31]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i18 (.D(SLO_buf[32]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i19 (.D(SLO_buf[33]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i20 (.D(SLO_buf[34]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i21 (.D(SLO_buf[35]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i22 (.D(SLO_buf[36]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i23 (.D(SLO_buf[37]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i24 (.D(SLO_buf[38]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i25 (.D(SLO_buf[39]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i26 (.D(SLO_buf[40]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i27 (.D(SLO_buf[41]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i28 (.D(SLO_buf[42]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i29 (.D(SLO_buf[43]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i30 (.D(SLO_buf[44]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i31 (.D(SLO_buf[45]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(spi_data_out_r_39__N_5448[32]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i33 (.D(spi_data_out_r_39__N_5448[33]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i33.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i34 (.D(spi_data_out_r_39__N_5448[34]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i34.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i35 (.D(spi_data_out_r_39__N_5448[35]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5197[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i35.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i36 (.D(SLO_buf[10]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i36.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i37 (.D(SLO_buf[11]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i37.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i38 (.D(SLO_buf[12]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i38.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i39 (.D(SLO_buf[13]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5197[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i39.GSR = "DISABLED";
    LUT4 mux_158_i1_3_lut (.A(SLO_buf[14]), .B(SLO_buf[4]), .C(n47), .Z(spi_data_out_r_39__N_5448[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i1_3_lut.init = 16'hcaca;
    FD1P3AX Cnt_NSL_1782__i1 (.D(n53[1]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782__i1.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1782__i2 (.D(n53[2]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782__i2.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1782__i3 (.D(n53[3]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782__i3.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1782__i4 (.D(n53[4]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782__i4.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1782__i5 (.D(n53[5]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782__i5.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1782__i6 (.D(n53[6]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782__i6.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1782__i7 (.D(n53[7]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782__i7.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1782__i8 (.D(n53[8]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782__i8.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1782__i9 (.D(n53[9]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782__i9.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1782__i10 (.D(n53[10]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782__i10.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1782__i11 (.D(n53[11]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1782__i11.GSR = "DISABLED";
    PFUMX MA_Temp_I_205 (.BLUT(n28589), .ALUT(n28590), .C0(n18592), .Z(MA_Temp_N_5516)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;
    LUT4 i23982_4_lut (.A(NSL), .B(n30079), .C(n18592), .D(n30002), 
         .Z(NSL_N_5529)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C+(D))))) */ ;
    defparam i23982_4_lut.init = 16'h3b37;
    LUT4 i14194_3_lut_4_lut (.A(n30184), .B(n30183), .C(resetn_c), .D(n18592), 
         .Z(clk_1MHz_enable_68)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i14194_3_lut_4_lut.init = 16'h70f0;
    CCU2D add_564_9 (.A0(Cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21959), 
          .S0(n153[7]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_9.INIT0 = 16'h5aaa;
    defparam add_564_9.INIT1 = 16'h0000;
    defparam add_564_9.INJECT1_0 = "NO";
    defparam add_564_9.INJECT1_1 = "NO";
    CCU2D add_564_7 (.A0(Cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21958), 
          .COUT(n21959), .S0(n153[5]), .S1(n153[6]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_7.INIT0 = 16'h5aaa;
    defparam add_564_7.INIT1 = 16'h5aaa;
    defparam add_564_7.INJECT1_0 = "NO";
    defparam add_564_7.INJECT1_1 = "NO";
    CCU2D add_564_5 (.A0(Cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21957), 
          .COUT(n21958), .S0(n153[3]), .S1(n153[4]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_5.INIT0 = 16'h5aaa;
    defparam add_564_5.INIT1 = 16'h5aaa;
    defparam add_564_5.INJECT1_0 = "NO";
    defparam add_564_5.INJECT1_1 = "NO";
    CCU2D add_564_3 (.A0(Cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21956), 
          .COUT(n21957), .S0(n153[1]), .S1(n153[2]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_3.INIT0 = 16'h5aaa;
    defparam add_564_3.INIT1 = 16'h5aaa;
    defparam add_564_3.INJECT1_0 = "NO";
    defparam add_564_3.INJECT1_1 = "NO";
    CCU2D add_564_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n21956), 
          .S1(n153[0]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_1.INIT0 = 16'hF000;
    defparam add_564_1.INIT1 = 16'h5555;
    defparam add_564_1.INJECT1_0 = "NO";
    defparam add_564_1.INJECT1_1 = "NO";
    LUT4 i23989_3_lut (.A(n25979), .B(n23916), .C(n30199), .Z(clk_enable_221)) /* synthesis lut_function=(!(A (B (C)))) */ ;
    defparam i23989_3_lut.init = 16'h7f7f;
    LUT4 i1_2_lut_adj_817 (.A(\quad_homing[0] ), .B(pin_io_c_44), .Z(n25893)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(74[8:17])
    defparam i1_2_lut_adj_817.init = 16'h8888;
    LUT4 i2429_2_lut_rep_779 (.A(mode[0]), .B(mode[1]), .Z(n30179)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2429_2_lut_rep_779.init = 16'h8888;
    LUT4 i24086_2_lut_3_lut (.A(mode[0]), .B(mode[1]), .C(mode[2]), .Z(ENC_O_N_5498)) /* synthesis lut_function=(!(A (B+(C))+!A (C))) */ ;
    defparam i24086_2_lut_3_lut.init = 16'h0707;
    LUT4 i1_3_lut_rep_780 (.A(mode[1]), .B(mode[2]), .C(mode[0]), .Z(n30180)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_3_lut_rep_780.init = 16'hfbfb;
    LUT4 i24081_2_lut_4_lut (.A(mode[1]), .B(mode[2]), .C(mode[0]), .D(TX_IN_N_6565), 
         .Z(n7163)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i24081_2_lut_4_lut.init = 16'h00fb;
    LUT4 i1_2_lut_4_lut (.A(mode[1]), .B(mode[2]), .C(mode[0]), .D(Cnt[5]), 
         .Z(n26301)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_4_lut.init = 16'hfffb;
    LUT4 i1_3_lut_rep_685_4_lut (.A(Cnt[2]), .B(Cnt[3]), .C(Cnt[0]), .D(n23598), 
         .Z(n30085)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(109[8:17])
    defparam i1_3_lut_rep_685_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut (.A(Cnt[2]), .B(Cnt[3]), .C(Cnt[1]), .D(Cnt[0]), 
         .Z(n18498)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(109[8:17])
    defparam i1_3_lut_4_lut.init = 16'hfeee;
    LUT4 i1_3_lut_rep_783 (.A(Cnt_NSL[9]), .B(Cnt_NSL[8]), .C(Cnt_NSL[7]), 
         .Z(n30183)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_rep_783.init = 16'hfefe;
    LUT4 i1_2_lut_rep_679_4_lut (.A(Cnt_NSL[9]), .B(Cnt_NSL[8]), .C(Cnt_NSL[7]), 
         .D(n30184), .Z(n30079)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_rep_679_4_lut.init = 16'hfe00;
    LUT4 i1_2_lut_rep_784 (.A(Cnt_NSL[11]), .B(Cnt_NSL[10]), .Z(n30184)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i1_2_lut_rep_784.init = 16'h8888;
    LUT4 i23946_2_lut_rep_630_3_lut_4_lut (.A(Cnt_NSL[11]), .B(Cnt_NSL[10]), 
         .C(resetn_c), .D(n30183), .Z(clk_1MHz_enable_20)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i23946_2_lut_rep_630_3_lut_4_lut.init = 16'h8f0f;
    LUT4 i24150_4_lut (.A(n30086), .B(n26387), .C(n30180), .D(mode[2]), 
         .Z(clk_enable_1103)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C)))) */ ;
    defparam i24150_4_lut.init = 16'h0545;
    LUT4 i1_4_lut_adj_818 (.A(mode[1]), .B(mode[0]), .C(Cnt[4]), .D(n4), 
         .Z(n26387)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_818.init = 16'h8880;
    LUT4 i19098_2_lut (.A(\uart_slot_en[1] ), .B(\uart_slot_en[2] ), .Z(n23722)) /* synthesis lut_function=(A (B)) */ ;
    defparam i19098_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_819 (.A(clk_enable_641), .B(EM_STOP), .C(n25699), 
         .D(n23916), .Z(clk_enable_36)) /* synthesis lut_function=(A+!((C (D))+!B)) */ ;
    defparam i1_4_lut_adj_819.init = 16'haeee;
    LUT4 mux_158_i2_3_lut (.A(SLO_buf[15]), .B(SLO_buf[5]), .C(n47), .Z(spi_data_out_r_39__N_5448[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i2_3_lut.init = 16'hcaca;
    LUT4 mux_158_i3_3_lut (.A(SLO_buf[16]), .B(SLO_buf[6]), .C(n47), .Z(spi_data_out_r_39__N_5448[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i3_3_lut.init = 16'hcaca;
    LUT4 mux_158_i4_3_lut (.A(SLO_buf[17]), .B(SLO_buf[7]), .C(n47), .Z(spi_data_out_r_39__N_5448[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i4_3_lut.init = 16'hcaca;
    LUT4 mux_158_i5_3_lut (.A(SLO_buf[18]), .B(SLO_buf[8]), .C(n47), .Z(spi_data_out_r_39__N_5448[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i5_3_lut.init = 16'hcaca;
    LUT4 mux_158_i6_3_lut (.A(SLO_buf[19]), .B(SLO_buf[9]), .C(n47), .Z(spi_data_out_r_39__N_5448[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i6_3_lut.init = 16'hcaca;
    LUT4 mux_158_i7_3_lut (.A(SLO_buf[20]), .B(SLO_buf[10]), .C(n47), 
         .Z(spi_data_out_r_39__N_5448[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i7_3_lut.init = 16'hcaca;
    LUT4 mux_158_i8_3_lut (.A(SLO_buf[21]), .B(SLO_buf[11]), .C(n47), 
         .Z(spi_data_out_r_39__N_5448[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i8_3_lut.init = 16'hcaca;
    LUT4 mux_158_i9_3_lut (.A(SLO_buf[22]), .B(SLO_buf[12]), .C(n47), 
         .Z(spi_data_out_r_39__N_5448[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i9_3_lut.init = 16'hcaca;
    LUT4 mux_158_i10_3_lut (.A(SLO_buf[23]), .B(SLO_buf[13]), .C(n47), 
         .Z(spi_data_out_r_39__N_5448[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i10_3_lut.init = 16'hcaca;
    LUT4 mux_158_i11_3_lut (.A(SLO_buf[24]), .B(SLO_buf[14]), .C(n47), 
         .Z(spi_data_out_r_39__N_5448[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i11_3_lut.init = 16'hcaca;
    LUT4 mux_158_i12_3_lut (.A(SLO_buf[25]), .B(SLO_buf[15]), .C(n47), 
         .Z(spi_data_out_r_39__N_5448[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i12_3_lut.init = 16'hcaca;
    LUT4 mux_158_i13_3_lut (.A(SLO_buf[26]), .B(SLO_buf[16]), .C(n47), 
         .Z(spi_data_out_r_39__N_5448[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i13_3_lut.init = 16'hcaca;
    LUT4 mux_158_i14_3_lut (.A(SLO_buf[27]), .B(SLO_buf[17]), .C(n47), 
         .Z(spi_data_out_r_39__N_5448[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i14_3_lut.init = 16'hcaca;
    LUT4 mux_158_i15_3_lut (.A(SLO_buf[28]), .B(SLO_buf[18]), .C(n47), 
         .Z(spi_data_out_r_39__N_5448[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i15_3_lut.init = 16'hcaca;
    LUT4 mux_158_i16_3_lut (.A(SLO_buf[29]), .B(SLO_buf[19]), .C(n47), 
         .Z(spi_data_out_r_39__N_5448[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i16_3_lut.init = 16'hcaca;
    LUT4 mux_158_i33_3_lut (.A(SLO_buf[6]), .B(SLO_buf[0]), .C(n47), .Z(spi_data_out_r_39__N_5448[32])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i33_3_lut.init = 16'hcaca;
    LUT4 mux_158_i34_3_lut (.A(SLO_buf[7]), .B(SLO_buf[1]), .C(n47), .Z(spi_data_out_r_39__N_5448[33])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i34_3_lut.init = 16'hcaca;
    LUT4 mux_158_i35_3_lut (.A(SLO_buf[8]), .B(SLO_buf[2]), .C(n47), .Z(spi_data_out_r_39__N_5448[34])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i35_3_lut.init = 16'hcaca;
    LUT4 mux_158_i36_3_lut (.A(SLO_buf[9]), .B(SLO_buf[3]), .C(n47), .Z(spi_data_out_r_39__N_5448[35])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i36_3_lut.init = 16'hcaca;
    LUT4 digital_output_r_I_0_547_3_lut (.A(digital_output_r), .B(UC_TXD0_c), 
         .C(OW_ID_N_5491), .Z(OW_ID_N_5490)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[16] 91[59])
    defparam digital_output_r_I_0_547_3_lut.init = 16'hcaca;
    LUT4 i4_4_lut (.A(n30207), .B(n30050), .C(n30120), .D(mode[0]), 
         .Z(OW_ID_N_5491)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i4_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_rep_807 (.A(mode[1]), .B(mode[2]), .Z(n30207)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i1_2_lut_rep_807.init = 16'heeee;
    LUT4 i2988_2_lut_3_lut_4_lut (.A(mode[1]), .B(mode[2]), .C(pin_io_out_49), 
         .D(mode[0]), .Z(\quad_b[4] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i2988_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i2987_2_lut_3_lut_4_lut (.A(mode[1]), .B(mode[2]), .C(pin_io_c_48), 
         .D(mode[0]), .Z(\quad_a[4] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i2987_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i24025_2_lut_3_lut_4_lut (.A(n30079), .B(resetn_c), .C(n18592), 
         .D(n18530), .Z(clk_1MHz_enable_8)) /* synthesis lut_function=(!(A (C (D))+!A (B+(C (D))))) */ ;
    defparam i24025_2_lut_3_lut_4_lut.init = 16'h0bbb;
    LUT4 i1_2_lut_3_lut (.A(Cnt[5]), .B(n30085), .C(Cnt[1]), .Z(n4)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(133[16:19])
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i23897_1_lut_2_lut_3_lut_4_lut (.A(Cnt[5]), .B(n30085), .C(MA_Temp), 
         .D(n30148), .Z(n28589)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(133[16:19])
    defparam i23897_1_lut_2_lut_3_lut_4_lut.init = 16'he1f0;
    LUT4 i23898_1_lut_4_lut (.A(MA_Temp), .B(n18530), .C(n28322), .D(n30085), 
         .Z(n28590)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A (B+((D)+!C)))) */ ;
    defparam i23898_1_lut_4_lut.init = 16'h2212;
    FD1P3IX SLO__i43 (.D(SLO[41]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i43.GSR = "DISABLED";
    FD1P3IX SLO__i44 (.D(SLO[42]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i44.GSR = "DISABLED";
    FD1P3IX SLO__i41 (.D(SLO[39]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i41.GSR = "DISABLED";
    FD1P3IX SLO__i45 (.D(SLO[43]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i45.GSR = "DISABLED";
    FD1P3IX SLO__i42 (.D(SLO[40]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i42.GSR = "DISABLED";
    FD1P3IX SLO__i46 (.D(SLO[44]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i46.GSR = "DISABLED";
    FD1P3IX SLO__i31 (.D(SLO[29]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i31.GSR = "DISABLED";
    FD1P3IX SLO__i35 (.D(SLO[33]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i35.GSR = "DISABLED";
    FD1P3IX SLO__i38 (.D(SLO[36]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i38.GSR = "DISABLED";
    FD1P3IX SLO__i32 (.D(SLO[30]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i32.GSR = "DISABLED";
    FD1P3IX SLO__i36 (.D(SLO[34]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i36.GSR = "DISABLED";
    FD1P3IX SLO__i39 (.D(SLO[37]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i39.GSR = "DISABLED";
    FD1P3IX SLO__i29 (.D(SLO[27]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i29.GSR = "DISABLED";
    FD1P3IX SLO__i33 (.D(SLO[31]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i33.GSR = "DISABLED";
    FD1P3IX SLO__i30 (.D(SLO[28]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i30.GSR = "DISABLED";
    FD1P3IX SLO__i34 (.D(SLO[32]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i34.GSR = "DISABLED";
    FD1P3IX SLO__i37 (.D(SLO[35]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i37.GSR = "DISABLED";
    FD1P3IX SLO__i40 (.D(SLO[38]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i40.GSR = "DISABLED";
    FD1P3IX SLO__i20 (.D(SLO[18]), .SP(clk_enable_1103), .CD(GND_net), 
            .CK(clk), .Q(SLO[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i20.GSR = "DISABLED";
    FD1P3IX SLO__i23 (.D(SLO[21]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i23.GSR = "DISABLED";
    FD1P3IX SLO__i26 (.D(SLO[24]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i26.GSR = "DISABLED";
    FD1P3IX SLO__i24 (.D(SLO[22]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i24.GSR = "DISABLED";
    FD1P3IX SLO__i27 (.D(SLO[25]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i27.GSR = "DISABLED";
    FD1P3IX SLO__i18 (.D(SLO[16]), .SP(clk_enable_1103), .CD(GND_net), 
            .CK(clk), .Q(SLO[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i18.GSR = "DISABLED";
    FD1P3IX SLO__i21 (.D(SLO[19]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i21.GSR = "DISABLED";
    FD1P3IX SLO__i19 (.D(SLO[17]), .SP(clk_enable_1103), .CD(GND_net), 
            .CK(clk), .Q(SLO[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i19.GSR = "DISABLED";
    FD1P3IX SLO__i22 (.D(SLO[20]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i22.GSR = "DISABLED";
    FD1P3IX SLO__i25 (.D(SLO[23]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i25.GSR = "DISABLED";
    FD1P3IX SLO__i28 (.D(SLO[26]), .SP(clk_enable_1103), .CD(n12496), 
            .CK(clk), .Q(SLO[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i28.GSR = "DISABLED";
    FD1P3IX SLO__i8 (.D(SLO[6]), .SP(clk_enable_1103), .CD(GND_net), .CK(clk), 
            .Q(SLO[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i8.GSR = "DISABLED";
    FD1P3IX SLO__i12 (.D(SLO[10]), .SP(clk_enable_1103), .CD(GND_net), 
            .CK(clk), .Q(SLO[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i12.GSR = "DISABLED";
    FD1P3IX SLO__i15 (.D(SLO[13]), .SP(clk_enable_1103), .CD(GND_net), 
            .CK(clk), .Q(SLO[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i15.GSR = "DISABLED";
    FD1P3IX SLO__i9 (.D(SLO[7]), .SP(clk_enable_1103), .CD(GND_net), .CK(clk), 
            .Q(SLO[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i9.GSR = "DISABLED";
    FD1P3IX SLO__i13 (.D(SLO[11]), .SP(clk_enable_1103), .CD(GND_net), 
            .CK(clk), .Q(SLO[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i13.GSR = "DISABLED";
    FD1P3IX SLO__i16 (.D(SLO[14]), .SP(clk_enable_1103), .CD(GND_net), 
            .CK(clk), .Q(SLO[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i16.GSR = "DISABLED";
    FD1P3IX SLO__i6 (.D(SLO[4]), .SP(clk_enable_1103), .CD(GND_net), .CK(clk), 
            .Q(SLO[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i6.GSR = "DISABLED";
    FD1P3IX SLO__i10 (.D(SLO[8]), .SP(clk_enable_1103), .CD(GND_net), 
            .CK(clk), .Q(SLO[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i10.GSR = "DISABLED";
    FD1P3IX SLO__i7 (.D(SLO[5]), .SP(clk_enable_1103), .CD(GND_net), .CK(clk), 
            .Q(SLO[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i7.GSR = "DISABLED";
    FD1P3IX SLO__i11 (.D(SLO[9]), .SP(clk_enable_1103), .CD(GND_net), 
            .CK(clk), .Q(SLO[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i11.GSR = "DISABLED";
    FD1P3IX SLO__i14 (.D(SLO[12]), .SP(clk_enable_1103), .CD(GND_net), 
            .CK(clk), .Q(SLO[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i14.GSR = "DISABLED";
    FD1P3IX SLO__i17 (.D(SLO[15]), .SP(clk_enable_1103), .CD(GND_net), 
            .CK(clk), .Q(SLO[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i17.GSR = "DISABLED";
    FD1P3IX SLO__i3 (.D(SLO[1]), .SP(clk_enable_1103), .CD(GND_net), .CK(clk), 
            .Q(SLO[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i3.GSR = "DISABLED";
    FD1P3IX SLO__i4 (.D(SLO[2]), .SP(clk_enable_1103), .CD(GND_net), .CK(clk), 
            .Q(SLO[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i4.GSR = "DISABLED";
    FD1P3AX NSL_484 (.D(NSL_N_5529), .SP(clk_1MHz_enable_68), .CK(clk_1MHz), 
            .Q(NSL)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam NSL_484.GSR = "DISABLED";
    FD1P3IX SLO__i2 (.D(SLO[0]), .SP(clk_enable_1103), .CD(GND_net), .CK(clk), 
            .Q(SLO[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i2.GSR = "DISABLED";
    FD1P3IX SLO__i5 (.D(SLO[3]), .SP(clk_enable_1103), .CD(GND_net), .CK(clk), 
            .Q(SLO[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i5.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_728 (.A(mode[2]), .B(mode[0]), .Z(n30128)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_rep_728.init = 16'heeee;
    LUT4 i2986_2_lut_3_lut_4_lut (.A(mode[2]), .B(mode[0]), .C(pin_io_c_44), 
         .D(mode[1]), .Z(\pin_intrpt[14] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2986_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_2_lut_rep_655_3_lut (.A(mode[2]), .B(mode[0]), .C(mode[1]), 
         .Z(n30055)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_rep_655_3_lut.init = 16'hfefe;
    LUT4 i24083_3_lut_4_lut (.A(mode[2]), .B(mode[0]), .C(mode[1]), .D(OW_ID_N_5491), 
         .Z(OW_ID_N_5496)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C+(D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i24083_3_lut_4_lut.init = 16'h00ef;
    LUT4 i2952_1_lut_2_lut_3_lut (.A(mode[2]), .B(mode[0]), .C(mode[1]), 
         .Z(n7266)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2952_1_lut_2_lut_3_lut.init = 16'h0101;
    LUT4 i2984_2_lut_3_lut_4_lut (.A(mode[2]), .B(mode[0]), .C(pin_io_c_42), 
         .D(mode[1]), .Z(\pin_intrpt[12] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2984_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2985_2_lut_3_lut_4_lut (.A(mode[2]), .B(mode[0]), .C(pin_io_c_43), 
         .D(mode[1]), .Z(\pin_intrpt[13] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2985_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i12977_2_lut_3_lut (.A(n18530), .B(n18592), .C(n153[0]), .Z(n199[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i12977_2_lut_3_lut.init = 16'h7070;
    LUT4 i13454_2_lut_3_lut (.A(n18530), .B(n18592), .C(n153[7]), .Z(n199[7])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13454_2_lut_3_lut.init = 16'h7070;
    LUT4 i13453_2_lut_3_lut (.A(n18530), .B(n18592), .C(n153[6]), .Z(n199[6])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13453_2_lut_3_lut.init = 16'h7070;
    LUT4 i13452_2_lut_3_lut (.A(n18530), .B(n18592), .C(n153[5]), .Z(n199[5])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13452_2_lut_3_lut.init = 16'h7070;
    LUT4 i13451_2_lut_3_lut (.A(n18530), .B(n18592), .C(n153[4]), .Z(n199[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13451_2_lut_3_lut.init = 16'h7070;
    LUT4 i23986_2_lut_rep_746 (.A(MA_Temp), .B(clk_1MHz), .Z(n30146)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i23986_2_lut_rep_746.init = 16'h7777;
    LUT4 i24158_2_lut_3_lut_4_lut (.A(MA_Temp), .B(clk_1MHz), .C(n30180), 
         .D(prev_MA), .Z(n12496)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i24158_2_lut_3_lut_4_lut.init = 16'h0007;
    LUT4 i13450_2_lut_3_lut (.A(n18530), .B(n18592), .C(n153[3]), .Z(n199[3])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13450_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_686_3_lut (.A(MA_Temp), .B(clk_1MHz), .C(prev_MA), 
         .Z(n30086)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i1_2_lut_rep_686_3_lut.init = 16'hf8f8;
    LUT4 i13449_2_lut_3_lut (.A(n18530), .B(n18592), .C(n153[2]), .Z(n199[2])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13449_2_lut_3_lut.init = 16'h7070;
    LUT4 i13158_2_lut_rep_748 (.A(Cnt[4]), .B(Cnt[1]), .Z(n30148)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13158_2_lut_rep_748.init = 16'h8888;
    LUT4 i13448_2_lut_3_lut (.A(n18530), .B(n18592), .C(n153[1]), .Z(n199[1])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13448_2_lut_3_lut.init = 16'h7070;
    LUT4 i23620_2_lut_3_lut (.A(Cnt[4]), .B(Cnt[1]), .C(Cnt[5]), .Z(n28322)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i23620_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_602_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(n30085), 
         .D(Cnt[5]), .Z(n30002)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_rep_602_3_lut_4_lut.init = 16'hfff7;
    
endmodule
//
// Verilog Description of module spi_slave_top
//

module spi_slave_top (spi_addr_r, clk, n30080, n30185, spi_data_valid_r, 
            spi_data_valid, n23916, n30035, \spi_data_r[0] , clk_enable_161, 
            spi_scsn_c, spi_addr_valid, spi_cmd_valid, \spi_data_r[31] , 
            \spi_data_r[30] , \spi_data_r[29] , \spi_data_r[28] , \spi_data_r[27] , 
            \spi_data_r[26] , \spi_data_r[25] , \spi_data_r[24] , \spi_data_r[23] , 
            \spi_data_r[22] , \spi_data_r[21] , \spi_data_r[20] , \spi_data_r[19] , 
            \spi_data_r[18] , \spi_data_r[17] , \spi_data_r[16] , spi_cmd_r, 
            n28328, n26327, \spi_data_r[15] , \spi_data_r[14] , \spi_data_r[13] , 
            \spi_data_r[12] , \spi_data_r[11] , \spi_data_r[10] , \spi_data_r[9] , 
            \spi_data_r[8] , \spi_data_r[7] , \spi_data_r[6] , \spi_data_r[5] , 
            \spi_data_r[4] , \spi_data_r[3] , \spi_data_r[2] , \spi_data_r[1] , 
            \spi_data_out_r[0] , n26621, n26819, n27013, n27015, n30144, 
            n30155, n18440, n28524, n4, n30044, n23526, n26545, 
            n30151, n30094, quad_set_valid_N_1158, n23732, n26497, 
            n30209, n28260, n30214, \spi_cmd[2] , \spi_data_out_r[1] , 
            \spi_data_out_r[3] , \spi_data_out_r[4] , \spi_data_out_r[5] , 
            \spi_data_out_r[6] , \spi_data_out_r[7] , \spi_data_out_r_39__N_5197[8] , 
            n16, spi_data_out_r_39__N_5237, \spi_data_out_r[10] , \spi_data_out_r[11] , 
            \spi_data_out_r[12] , \spi_data_out_r[13] , \spi_data_out_r[14] , 
            \spi_data_out_r[15] , \spi_data_out_r[16] , \spi_data_out_r[17] , 
            \spi_data_out_r[18] , \spi_data_out_r[19] , \spi_data_out_r[20] , 
            \spi_data_out_r[21] , \spi_data_out_r[22] , \spi_data_out_r[23] , 
            \spi_data_out_r[24] , \spi_data_out_r[25] , \spi_data_out_r[26] , 
            \spi_data_out_r[27] , \spi_data_out_r[28] , \spi_data_out_r[29] , 
            \spi_data_out_r[30] , \spi_data_out_r[31] , \spi_data_out_r[32] , 
            \spi_data_out_r[33] , \spi_data_out_r[34] , \spi_data_out_r[35] , 
            \spi_data_out_r[36] , \spi_data_out_r[37] , \spi_data_out_r[38] , 
            \spi_data_out_r[39] , \spi_data_out_r_39__N_5540[8] , n18, 
            spi_data_out_r_39__N_5580, \spi_data_out_r_39__N_4168[8] , n3, 
            spi_data_out_r_39__N_4208, \spi_data_out_r_39__N_5883[8] , \spi_data_out_r_39__N_4854[8] , 
            spi_data_out_r_39__N_5923, spi_data_out_r_39__N_4894, \spi_data_out_r_39__N_2109[8] , 
            n5, spi_data_out_r_39__N_2149, \spi_data_out_r_39__N_1404[8] , 
            \spi_data_out_r_39__N_934[8] , spi_data_out_r_39__N_1444, spi_data_out_r_39__N_974, 
            n28384, \spi_data_out_r_39__N_2344[8] , \spi_data_out_r_39__N_1874[8] , 
            spi_data_out_r_39__N_2384, spi_data_out_r_39__N_1914, \spi_data_out_r_39__N_4168[9] , 
            n16_adj_329, \spi_data_out_r_39__N_5883[9] , n21, \spi_data_out_r_39__N_4854[9] , 
            n2, \spi_data_out_r_39__N_5197[9] , \spi_data_out_r_39__N_4511[9] , 
            spi_data_out_r_39__N_4551, \spi_data_out_r_39__N_1874[9] , n5_adj_330, 
            \spi_data_out_r_39__N_2344[9] , \spi_data_out_r_39__N_2109[9] , 
            \spi_data_out_r_39__N_1404[9] , \spi_data_out_r_39__N_1169[9] , 
            spi_data_out_r_39__N_1209, n21_adj_331, n19, \spi_data_out_r_39__N_5197[2] , 
            n22, \spi_data_out_r_39__N_2863[2] , \spi_data_out_r_39__N_2721[2] , 
            clear_intrpt, clear_intrpt_adj_332, \spi_data_out_r_39__N_4511[2] , 
            \spi_data_out_r_39__N_4168[2] , \spi_data_out_r_39__N_3005[2] , 
            n14, n9, clear_intrpt_adj_333, \spi_data_out_r_39__N_2792[2] , 
            \spi_data_out_r_39__N_2650[2] , clear_intrpt_adj_334, clear_intrpt_adj_335, 
            \spi_data_out_r_39__N_1169[2] , n7, \spi_data_out_r_39__N_1639[2] , 
            \spi_data_out_r_39__N_1404[2] , spi_data_out_r_39__N_1679, \spi_data_out_r_39__N_1874[2] , 
            \spi_data_out_r_39__N_2344[2] , \spi_data_out_r_39__N_3825[2] , 
            \spi_data_out_r_39__N_934[2] , spi_data_out_r_39__N_3865, n25721, 
            n28358, n26435, n26521, n30090, n26569, n24066, n28340, 
            quad_set_valid_N_1393, n30071, n25571, n26243, n30062, 
            n25859, resetn_c, n30210, n30213, n30023, n29995, n29996, 
            clk_enable_254, clk_enable_259, n30070, n29993, n25643, 
            n30064, n23537, n31069, GND_net, spi_mosi_oe, spi_mosi_o, 
            spi_miso_oe, spi_miso_o, spi_clk_oe, spi_clk_o, spi_mosi_i, 
            spi_miso_i, spi_clk_i, VCC_net, quad_buffer, quad_count, 
            \spi_data_out_r_39__N_1083[31] , \spi_data_out_r_39__N_1083[29] , 
            \spi_data_out_r_39__N_1083[19] , \spi_data_out_r_39__N_1083[18] , 
            quad_buffer_adj_644, quad_count_adj_645, \spi_data_out_r_39__N_2023[26] , 
            n30198, n32, clear_intrpt_N_2717, n47, clear_intrpt_N_2930, 
            clear_intrpt_N_2788, clear_intrpt_N_2859, n47_adj_400, quad_buffer_adj_646, 
            quad_count_adj_647, \spi_data_out_r_39__N_2493[29] , \spi_data_out_r_39__N_2493[28] , 
            \spi_data_out_r_39__N_2493[27] , \spi_data_out_r_39__N_2493[26] , 
            n29997, n29991, \spi_data_out_r_39__N_2493[25] , \spi_data_out_r_39__N_2493[24] , 
            \spi_data_out_r_39__N_2493[23] , \spi_data_out_r_39__N_2493[22] , 
            \spi_data_out_r_39__N_2493[21] , \spi_data_out_r_39__N_2493[20] , 
            \spi_data_out_r_39__N_2493[19] , \spi_data_out_r_39__N_2493[18] , 
            \spi_data_out_r_39__N_2493[17] , \spi_data_out_r_39__N_2493[16] , 
            \spi_data_out_r_39__N_2493[15] , \spi_data_out_r_39__N_2493[14] , 
            \spi_data_out_r_39__N_2493[13] , \spi_data_out_r_39__N_2493[12] , 
            \spi_data_out_r_39__N_2493[11] , \spi_data_out_r_39__N_2493[10] , 
            \spi_data_out_r_39__N_2493[9] , \spi_data_out_r_39__N_2493[8] , 
            \spi_data_out_r_39__N_2493[7] , \spi_data_out_r_39__N_1083[9] , 
            \spi_data_out_r_39__N_1083[8] , \spi_data_out_r_39__N_2493[6] , 
            \spi_data_out_r_39__N_2493[5] , \spi_data_out_r_39__N_2493[4] , 
            \spi_data_out_r_39__N_2493[3] , \spi_data_out_r_39__N_2493[2] , 
            \spi_data_out_r_39__N_2493[1] , \spi_data_out_r_39__N_2023[20] , 
            quad_buffer_adj_648, quad_count_adj_649, \spi_data_out_r_39__N_2258[0] , 
            \spi_data_out_r_39__N_2258[31] , \spi_data_out_r_39__N_2258[30] , 
            \spi_data_out_r_39__N_2258[29] , \spi_data_out_r_39__N_2258[28] , 
            \spi_data_out_r_39__N_2258[27] , \spi_data_out_r_39__N_2258[26] , 
            n26779, \spi_data_out_r_39__N_2258[25] , \spi_data_out_r_39__N_2258[24] , 
            \spi_data_out_r_39__N_1083[22] , \spi_data_out_r_39__N_2258[23] , 
            \spi_data_out_r_39__N_2258[22] , \spi_data_out_r_39__N_2258[21] , 
            \spi_data_out_r_39__N_2258[20] , \spi_data_out_r_39__N_2258[19] , 
            \spi_data_out_r_39__N_2258[18] , n47_adj_529, \spi_data_out_r_39__N_2258[17] , 
            \spi_data_out_r_39__N_2258[16] , \spi_data_out_r_39__N_2258[15] , 
            \spi_data_out_r_39__N_2258[14] , \spi_data_out_r_39__N_2258[13] , 
            \spi_data_out_r_39__N_2258[12] , \spi_data_out_r_39__N_2258[11] , 
            \spi_data_out_r_39__N_2258[10] , \spi_data_out_r_39__N_2258[9] , 
            n30019, n47_adj_530, \spi_data_out_r_39__N_2258[8] , \spi_data_out_r_39__N_2258[7] , 
            n30027, n47_adj_531, \spi_data_out_r_39__N_2258[6] , \spi_data_out_r_39__N_2258[5] , 
            \spi_data_out_r_39__N_2258[4] , \spi_data_out_r_39__N_2258[3] , 
            \spi_data_out_r_39__N_1083[17] , \spi_data_out_r_39__N_2258[2] , 
            \spi_data_out_r_39__N_2023[19] , \spi_data_out_r_39__N_2258[1] , 
            \SLO_buf[4] , \SLO_buf[14] , \spi_data_out_r_39__N_5105[0] , 
            \SLO_buf[3] , \SLO_buf[9] , \spi_data_out_r_39__N_5105[35] , 
            \SLO_buf[2] , \SLO_buf[8] , \spi_data_out_r_39__N_5105[34] , 
            \SLO_buf[1] , \SLO_buf[7] , \spi_data_out_r_39__N_5105[33] , 
            quad_buffer_adj_650, quad_count_adj_651, \spi_data_out_r_39__N_1553[0] , 
            \spi_data_out_r_39__N_1553[31] , \SLO_buf[0] , \SLO_buf[6] , 
            \spi_data_out_r_39__N_5105[32] , \SLO_buf[19] , \SLO_buf[29] , 
            \spi_data_out_r_39__N_5105[15] , \spi_data_out_r_39__N_1553[30] , 
            \spi_data_out_r_39__N_1553[29] , \spi_data_out_r_39__N_1553[28] , 
            \spi_data_out_r_39__N_1553[27] , \SLO_buf[18] , \SLO_buf[28] , 
            \spi_data_out_r_39__N_5105[14] , \spi_data_out_r_39__N_1553[26] , 
            \SLO_buf[17] , \SLO_buf[27] , \spi_data_out_r_39__N_5105[13] , 
            \spi_data_out_r_39__N_2023[25] , \spi_data_out_r_39__N_1553[25] , 
            \spi_data_out_r_39__N_1553[24] , \SLO_buf[16] , \SLO_buf[26] , 
            \spi_data_out_r_39__N_5105[12] , \spi_data_out_r_39__N_1553[23] , 
            \SLO_buf[15] , \SLO_buf[25] , \spi_data_out_r_39__N_5105[11] , 
            \SLO_buf[24] , \spi_data_out_r_39__N_5105[10] , \spi_data_out_r_39__N_1553[22] , 
            \SLO_buf[13] , \SLO_buf[23] , \spi_data_out_r_39__N_5105[9] , 
            \spi_data_out_r_39__N_1553[21] , \spi_data_out_r_39__N_1553[20] , 
            \spi_data_out_r_39__N_1553[19] , \spi_data_out_r_39__N_1553[18] , 
            \spi_data_out_r_39__N_1553[17] , \spi_data_out_r_39__N_1553[16] , 
            \spi_data_out_r_39__N_1083[16] , \spi_data_out_r_39__N_1553[15] , 
            \spi_data_out_r_39__N_1553[14] , \spi_data_out_r_39__N_1553[13] , 
            \spi_data_out_r_39__N_1083[15] , \SLO_buf[12] , \SLO_buf[22] , 
            \spi_data_out_r_39__N_5105[8] , \spi_data_out_r_39__N_1553[12] , 
            \SLO_buf[11] , \SLO_buf[21] , \spi_data_out_r_39__N_5105[7] , 
            \spi_data_out_r_39__N_1553[11] , \SLO_buf[10] , \SLO_buf[20] , 
            \spi_data_out_r_39__N_5105[6] , \spi_data_out_r_39__N_5105[5] , 
            \spi_data_out_r_39__N_1553[10] , \spi_data_out_r_39__N_5105[4] , 
            \spi_data_out_r_39__N_1553[9] , \spi_data_out_r_39__N_1553[8] , 
            \spi_data_out_r_39__N_1553[7] , \spi_data_out_r_39__N_1553[6] , 
            \spi_data_out_r_39__N_5105[3] , \spi_data_out_r_39__N_1553[5] , 
            \spi_data_out_r_39__N_1553[4] , \spi_data_out_r_39__N_1553[3] , 
            \spi_data_out_r_39__N_2023[18] , \spi_data_out_r_39__N_1553[2] , 
            \spi_data_out_r_39__N_1553[1] , n47_adj_596, \spi_data_out_r_39__N_5105[2] , 
            \SLO_buf[5] , \spi_data_out_r_39__N_5105[1] , spi_data_out_r_39__N_2338, 
            n47_adj_597, \spi_data_out_r_39__N_1083[14] , \spi_data_out_r_39__N_1083[13] , 
            n30102, \SLO_buf[4]_adj_598 , \SLO_buf[14]_adj_599 , \spi_data_out_r_39__N_4419[0] , 
            \SLO_buf[3]_adj_600 , \SLO_buf[9]_adj_601 , \spi_data_out_r_39__N_4419[35] , 
            spi_data_out_r_39__N_4505, \spi_data_out_r_39__N_2023[17] , 
            \spi_data_out_r_39__N_2023[16] , \spi_data_out_r_39__N_1083[7] , 
            \spi_data_out_r_39__N_1083[6] , \spi_data_out_r_39__N_1083[20] , 
            \spi_data_out_r_39__N_2023[15] , \status_cntr[12] , n25212, 
            \SLO_buf[2]_adj_602 , \SLO_buf[8]_adj_603 , \spi_data_out_r_39__N_4419[34] , 
            \spi_data_out_r_39__N_2023[14] , \SLO_buf[1]_adj_604 , \SLO_buf[7]_adj_605 , 
            \spi_data_out_r_39__N_4419[33] , \SLO_buf[0]_adj_606 , \SLO_buf[6]_adj_607 , 
            \spi_data_out_r_39__N_4419[32] , clear_intrpt_N_3072, \spi_data_out_r_39__N_2023[13] , 
            \SLO_buf[19]_adj_608 , \SLO_buf[29]_adj_609 , \spi_data_out_r_39__N_4419[15] , 
            \spi_data_out_r_39__N_1083[5] , \spi_data_out_r_39__N_1083[4] , 
            \spi_data_out_r_39__N_2023[12] , \SLO_buf[18]_adj_610 , \SLO_buf[28]_adj_611 , 
            \spi_data_out_r_39__N_4419[14] , \SLO_buf[17]_adj_612 , \SLO_buf[27]_adj_613 , 
            \spi_data_out_r_39__N_4419[13] , \spi_data_out_r_39__N_1083[12] , 
            spi_data_out_r_39__N_4848, \spi_data_out_r_39__N_1083[3] , \spi_data_out_r_39__N_1083[2] , 
            \spi_data_out_r_39__N_2023[11] , \SLO_buf[16]_adj_614 , \SLO_buf[26]_adj_615 , 
            \spi_data_out_r_39__N_4419[12] , \spi_data_out_r_39__N_2023[10] , 
            \SLO_buf[15]_adj_616 , \SLO_buf[25]_adj_617 , \spi_data_out_r_39__N_4419[11] , 
            \SLO_buf[24]_adj_618 , \spi_data_out_r_39__N_4419[10] , \SLO_buf[13]_adj_619 , 
            \SLO_buf[23]_adj_620 , \spi_data_out_r_39__N_4419[9] , \SLO_buf[12]_adj_621 , 
            \SLO_buf[22]_adj_622 , \spi_data_out_r_39__N_4419[8] , n25885, 
            n30087, \quad_homing[1] , n1, clk_enable_686, clk_enable_260, 
            clear_intrpt_adj_623, intrpt_out_N_2642, intrpt_out_N_3068, 
            clk_enable_263, clk_enable_807, n12467, n20647, n18654, 
            n12435, n26873, clk_enable_320, n25877, n30075, \quad_homing[1]_adj_624 , 
            n1_adj_625, n30199, n26821, clk_enable_684, n26089, n26091, 
            clk_enable_255, EM_STOP, clk_enable_23, n26947, clk_enable_253, 
            pwm_out_N_3169, pwm_out_N_3153, clk_enable_15, n26107, n26113, 
            clear_intrpt_adj_626, intrpt_out_N_2997, clk_enable_687, n30045, 
            clk_enable_759, clk_enable_727, n11008, pwm_out_1_N_6491, 
            clk_enable_613, n26957, clk_enable_520, clk_enable_232, 
            clk_enable_28, clk_enable_226, clk_enable_639, pwm_out_3_N_6530, 
            clk_enable_1105, pwm_out_4_N_6549, clk_enable_1107, clk_enable_757, 
            clk_enable_245, pwm_out_2_N_6511, clk_enable_22, clk_enable_488, 
            n26633, clk_enable_641, clk_enable_638, clk_enable_959, 
            clk_enable_235, intrpt_out_N_2713, n57, reset_r_N_4129, 
            clk_enable_761, n29998, clk_enable_738, n25881, n30095, 
            \quad_homing[1]_adj_627 , n1_adj_628, clk_enable_652, quad_set_valid_N_2098, 
            clk_enable_683, clk_enable_211, n2109, n25893, n30055, 
            \quad_homing[1]_adj_629 , n1_adj_630, n25869, n30043, \quad_homing[1]_adj_631 , 
            n1_adj_632, n25873, n30091, \quad_homing[1]_adj_633 , n1_adj_634, 
            n28476, clk_enable_32, intrpt_out_N_2855, clk_enable_178, 
            intrpt_out_N_2784, clk_enable_842, clk_enable_627, clk_enable_234, 
            quad_set_valid_N_2333, clk_enable_315, \SLO_buf[11]_adj_635 , 
            \SLO_buf[21]_adj_636 , \spi_data_out_r_39__N_4419[7] , clk_enable_256, 
            n29999, clk_enable_12, clk_enable_749, clk_enable_388, n26207, 
            clk_enable_898, clk_enable_180, n18_adj_637, n2193, \SLO_buf[10]_adj_638 , 
            \SLO_buf[20]_adj_639 , \spi_data_out_r_39__N_4419[6] , clk_enable_244, 
            intrpt_out_N_2926, pwm_out_1_N_6306, clk_100k_enable_1, n25889, 
            n30083, \quad_homing[1]_adj_640 , n1_adj_641, clk_enable_595, 
            n30039, \spi_data_out_r_39__N_2023[9] , \spi_data_out_r_39__N_1083[24] , 
            clear_intrpt_N_3001, \spi_data_out_r_39__N_2023[8] , \spi_data_out_r_39__N_1083[11] , 
            \spi_data_out_r_39__N_2023[7] , \spi_data_out_r_39__N_1083[27] , 
            \spi_data_out_r_39__N_4419[5] , \spi_data_out_r_39__N_4419[4] , 
            \spi_data_out_r_39__N_2023[6] , n27095, spi_data_out_r_39__N_1868, 
            n29992, \spi_data_out_r_39__N_4419[3] , \spi_data_out_r_39__N_2023[5] , 
            \spi_data_out_r_39__N_2023[24] , \spi_data_out_r_39__N_4419[2] , 
            spi_data_out_r_39__N_5191, spi_data_out_r_39__N_5534, spi_data_out_r_39__N_5877, 
            \spi_data_out_r_39__N_1083[23] , spi_data_out_r_39__N_6220, 
            \spi_data_out_r_39__N_2023[4] , \spi_data_out_r_39__N_2023[23] , 
            \spi_data_out_r_39__N_1083[1] , \spi_data_out_r_39__N_1083[26] , 
            spi_data_out_r_39__N_1398, \spi_data_out_r_39__N_1083[25] , 
            \spi_data_out_r_39__N_1083[30] , n30013, \spi_data_out_r_39__N_2023[3] , 
            \SLO_buf[5]_adj_642 , \spi_data_out_r_39__N_4419[1] , \spi_data_out_r_39__N_2023[2] , 
            \spi_data_out_r_39__N_2023[1] , \spi_data_out_r_39__N_1083[10] , 
            \spi_data_out_r_39__N_2023[0] , \spi_data_out_r_39__N_2023[22] , 
            n30007, clk_enable_38, \spi_data_out_r_39__N_2023[21] , n30020, 
            \spi_data_out_r_39__N_2023[31] , clk_enable_227, \spi_data_out_r_39__N_2023[30] , 
            \spi_data_out_r_39__N_2023[29] , \spi_data_out_r_39__N_1083[28] , 
            \spi_data_out_r_39__N_2023[28] , \spi_data_out_r_39__N_2023[27] , 
            \spi_data_out_r_39__N_1083[21] , n22554, pwm, n4_adj_643, 
            \status_cntr[11] , \spi_data_out_r_39__N_1083[0] , spi_data_out_r_39__N_2103, 
            spi_data_out_r_39__N_1163, \spi_data_out_r_39__N_2493[0] , \spi_data_out_r_39__N_2493[31] , 
            \spi_data_out_r_39__N_2493[30] , spi_data_out_r_39__N_1633, 
            spi_data_out_r_39__N_2573) /* synthesis syn_module_defined=1 */ ;
    output [7:0]spi_addr_r;
    input clk;
    output n30080;
    output n30185;
    output spi_data_valid_r;
    output spi_data_valid;
    input n23916;
    output n30035;
    output \spi_data_r[0] ;
    input clk_enable_161;
    input spi_scsn_c;
    output spi_addr_valid;
    output spi_cmd_valid;
    output \spi_data_r[31] ;
    output \spi_data_r[30] ;
    output \spi_data_r[29] ;
    output \spi_data_r[28] ;
    output \spi_data_r[27] ;
    output \spi_data_r[26] ;
    output \spi_data_r[25] ;
    output \spi_data_r[24] ;
    output \spi_data_r[23] ;
    output \spi_data_r[22] ;
    output \spi_data_r[21] ;
    output \spi_data_r[20] ;
    output \spi_data_r[19] ;
    output \spi_data_r[18] ;
    output \spi_data_r[17] ;
    output \spi_data_r[16] ;
    output [15:0]spi_cmd_r;
    input n28328;
    output n26327;
    output \spi_data_r[15] ;
    output \spi_data_r[14] ;
    output \spi_data_r[13] ;
    output \spi_data_r[12] ;
    output \spi_data_r[11] ;
    output \spi_data_r[10] ;
    output \spi_data_r[9] ;
    output \spi_data_r[8] ;
    output \spi_data_r[7] ;
    output \spi_data_r[6] ;
    output \spi_data_r[5] ;
    output \spi_data_r[4] ;
    output \spi_data_r[3] ;
    output \spi_data_r[2] ;
    output \spi_data_r[1] ;
    input \spi_data_out_r[0] ;
    input n26621;
    output n26819;
    input n27013;
    output n27015;
    output n30144;
    input n30155;
    input n18440;
    output n28524;
    input n4;
    output n30044;
    output n23526;
    input n26545;
    input n30151;
    input n30094;
    output quad_set_valid_N_1158;
    input n23732;
    input n26497;
    output n30209;
    input n28260;
    input n30214;
    output \spi_cmd[2] ;
    input \spi_data_out_r[1] ;
    input \spi_data_out_r[3] ;
    input \spi_data_out_r[4] ;
    input \spi_data_out_r[5] ;
    input \spi_data_out_r[6] ;
    input \spi_data_out_r[7] ;
    input \spi_data_out_r_39__N_5197[8] ;
    input n16;
    input spi_data_out_r_39__N_5237;
    input \spi_data_out_r[10] ;
    input \spi_data_out_r[11] ;
    input \spi_data_out_r[12] ;
    input \spi_data_out_r[13] ;
    input \spi_data_out_r[14] ;
    input \spi_data_out_r[15] ;
    input \spi_data_out_r[16] ;
    input \spi_data_out_r[17] ;
    input \spi_data_out_r[18] ;
    input \spi_data_out_r[19] ;
    input \spi_data_out_r[20] ;
    input \spi_data_out_r[21] ;
    input \spi_data_out_r[22] ;
    input \spi_data_out_r[23] ;
    input \spi_data_out_r[24] ;
    input \spi_data_out_r[25] ;
    input \spi_data_out_r[26] ;
    input \spi_data_out_r[27] ;
    input \spi_data_out_r[28] ;
    input \spi_data_out_r[29] ;
    input \spi_data_out_r[30] ;
    input \spi_data_out_r[31] ;
    input \spi_data_out_r[32] ;
    input \spi_data_out_r[33] ;
    input \spi_data_out_r[34] ;
    input \spi_data_out_r[35] ;
    input \spi_data_out_r[36] ;
    input \spi_data_out_r[37] ;
    input \spi_data_out_r[38] ;
    input \spi_data_out_r[39] ;
    input \spi_data_out_r_39__N_5540[8] ;
    input n18;
    input spi_data_out_r_39__N_5580;
    input \spi_data_out_r_39__N_4168[8] ;
    input n3;
    input spi_data_out_r_39__N_4208;
    input \spi_data_out_r_39__N_5883[8] ;
    input \spi_data_out_r_39__N_4854[8] ;
    input spi_data_out_r_39__N_5923;
    input spi_data_out_r_39__N_4894;
    input \spi_data_out_r_39__N_2109[8] ;
    input n5;
    input spi_data_out_r_39__N_2149;
    input \spi_data_out_r_39__N_1404[8] ;
    input \spi_data_out_r_39__N_934[8] ;
    input spi_data_out_r_39__N_1444;
    input spi_data_out_r_39__N_974;
    output n28384;
    input \spi_data_out_r_39__N_2344[8] ;
    input \spi_data_out_r_39__N_1874[8] ;
    input spi_data_out_r_39__N_2384;
    input spi_data_out_r_39__N_1914;
    input \spi_data_out_r_39__N_4168[9] ;
    input n16_adj_329;
    input \spi_data_out_r_39__N_5883[9] ;
    input n21;
    input \spi_data_out_r_39__N_4854[9] ;
    input n2;
    input \spi_data_out_r_39__N_5197[9] ;
    input \spi_data_out_r_39__N_4511[9] ;
    input spi_data_out_r_39__N_4551;
    input \spi_data_out_r_39__N_1874[9] ;
    input n5_adj_330;
    input \spi_data_out_r_39__N_2344[9] ;
    input \spi_data_out_r_39__N_2109[9] ;
    input \spi_data_out_r_39__N_1404[9] ;
    input \spi_data_out_r_39__N_1169[9] ;
    input spi_data_out_r_39__N_1209;
    input n21_adj_331;
    input n19;
    input \spi_data_out_r_39__N_5197[2] ;
    input n22;
    input \spi_data_out_r_39__N_2863[2] ;
    input \spi_data_out_r_39__N_2721[2] ;
    input clear_intrpt;
    input clear_intrpt_adj_332;
    input \spi_data_out_r_39__N_4511[2] ;
    input \spi_data_out_r_39__N_4168[2] ;
    input \spi_data_out_r_39__N_3005[2] ;
    input n14;
    input n9;
    input clear_intrpt_adj_333;
    input \spi_data_out_r_39__N_2792[2] ;
    input \spi_data_out_r_39__N_2650[2] ;
    input clear_intrpt_adj_334;
    input clear_intrpt_adj_335;
    input \spi_data_out_r_39__N_1169[2] ;
    input n7;
    input \spi_data_out_r_39__N_1639[2] ;
    input \spi_data_out_r_39__N_1404[2] ;
    input spi_data_out_r_39__N_1679;
    input \spi_data_out_r_39__N_1874[2] ;
    input \spi_data_out_r_39__N_2344[2] ;
    input \spi_data_out_r_39__N_3825[2] ;
    input \spi_data_out_r_39__N_934[2] ;
    input spi_data_out_r_39__N_3865;
    output n25721;
    input n28358;
    output n26435;
    input n26521;
    input n30090;
    input n26569;
    output n24066;
    input n28340;
    output quad_set_valid_N_1393;
    input n30071;
    output n25571;
    input n26243;
    input n30062;
    output n25859;
    input resetn_c;
    output n30210;
    output n30213;
    input n30023;
    output n29995;
    output n29996;
    output clk_enable_254;
    output clk_enable_259;
    output n30070;
    output n29993;
    output n25643;
    output n30064;
    output n23537;
    input n31069;
    input GND_net;
    output spi_mosi_oe;
    output spi_mosi_o;
    output spi_miso_oe;
    output spi_miso_o;
    output spi_clk_oe;
    output spi_clk_o;
    input spi_mosi_i;
    input spi_miso_i;
    input spi_clk_i;
    input VCC_net;
    input [31:0]quad_buffer;
    input [31:0]quad_count;
    output \spi_data_out_r_39__N_1083[31] ;
    output \spi_data_out_r_39__N_1083[29] ;
    output \spi_data_out_r_39__N_1083[19] ;
    output \spi_data_out_r_39__N_1083[18] ;
    input [31:0]quad_buffer_adj_644;
    input [31:0]quad_count_adj_645;
    output \spi_data_out_r_39__N_2023[26] ;
    output n30198;
    output n32;
    output clear_intrpt_N_2717;
    output n47;
    output clear_intrpt_N_2930;
    output clear_intrpt_N_2788;
    output clear_intrpt_N_2859;
    output n47_adj_400;
    input [31:0]quad_buffer_adj_646;
    input [31:0]quad_count_adj_647;
    output \spi_data_out_r_39__N_2493[29] ;
    output \spi_data_out_r_39__N_2493[28] ;
    output \spi_data_out_r_39__N_2493[27] ;
    output \spi_data_out_r_39__N_2493[26] ;
    output n29997;
    output n29991;
    output \spi_data_out_r_39__N_2493[25] ;
    output \spi_data_out_r_39__N_2493[24] ;
    output \spi_data_out_r_39__N_2493[23] ;
    output \spi_data_out_r_39__N_2493[22] ;
    output \spi_data_out_r_39__N_2493[21] ;
    output \spi_data_out_r_39__N_2493[20] ;
    output \spi_data_out_r_39__N_2493[19] ;
    output \spi_data_out_r_39__N_2493[18] ;
    output \spi_data_out_r_39__N_2493[17] ;
    output \spi_data_out_r_39__N_2493[16] ;
    output \spi_data_out_r_39__N_2493[15] ;
    output \spi_data_out_r_39__N_2493[14] ;
    output \spi_data_out_r_39__N_2493[13] ;
    output \spi_data_out_r_39__N_2493[12] ;
    output \spi_data_out_r_39__N_2493[11] ;
    output \spi_data_out_r_39__N_2493[10] ;
    output \spi_data_out_r_39__N_2493[9] ;
    output \spi_data_out_r_39__N_2493[8] ;
    output \spi_data_out_r_39__N_2493[7] ;
    output \spi_data_out_r_39__N_1083[9] ;
    output \spi_data_out_r_39__N_1083[8] ;
    output \spi_data_out_r_39__N_2493[6] ;
    output \spi_data_out_r_39__N_2493[5] ;
    output \spi_data_out_r_39__N_2493[4] ;
    output \spi_data_out_r_39__N_2493[3] ;
    output \spi_data_out_r_39__N_2493[2] ;
    output \spi_data_out_r_39__N_2493[1] ;
    output \spi_data_out_r_39__N_2023[20] ;
    input [31:0]quad_buffer_adj_648;
    input [31:0]quad_count_adj_649;
    output \spi_data_out_r_39__N_2258[0] ;
    output \spi_data_out_r_39__N_2258[31] ;
    output \spi_data_out_r_39__N_2258[30] ;
    output \spi_data_out_r_39__N_2258[29] ;
    output \spi_data_out_r_39__N_2258[28] ;
    output \spi_data_out_r_39__N_2258[27] ;
    output \spi_data_out_r_39__N_2258[26] ;
    output n26779;
    output \spi_data_out_r_39__N_2258[25] ;
    output \spi_data_out_r_39__N_2258[24] ;
    output \spi_data_out_r_39__N_1083[22] ;
    output \spi_data_out_r_39__N_2258[23] ;
    output \spi_data_out_r_39__N_2258[22] ;
    output \spi_data_out_r_39__N_2258[21] ;
    output \spi_data_out_r_39__N_2258[20] ;
    output \spi_data_out_r_39__N_2258[19] ;
    output \spi_data_out_r_39__N_2258[18] ;
    output n47_adj_529;
    output \spi_data_out_r_39__N_2258[17] ;
    output \spi_data_out_r_39__N_2258[16] ;
    output \spi_data_out_r_39__N_2258[15] ;
    output \spi_data_out_r_39__N_2258[14] ;
    output \spi_data_out_r_39__N_2258[13] ;
    output \spi_data_out_r_39__N_2258[12] ;
    output \spi_data_out_r_39__N_2258[11] ;
    output \spi_data_out_r_39__N_2258[10] ;
    output \spi_data_out_r_39__N_2258[9] ;
    output n30019;
    output n47_adj_530;
    output \spi_data_out_r_39__N_2258[8] ;
    output \spi_data_out_r_39__N_2258[7] ;
    output n30027;
    output n47_adj_531;
    output \spi_data_out_r_39__N_2258[6] ;
    output \spi_data_out_r_39__N_2258[5] ;
    output \spi_data_out_r_39__N_2258[4] ;
    output \spi_data_out_r_39__N_2258[3] ;
    output \spi_data_out_r_39__N_1083[17] ;
    output \spi_data_out_r_39__N_2258[2] ;
    output \spi_data_out_r_39__N_2023[19] ;
    output \spi_data_out_r_39__N_2258[1] ;
    input \SLO_buf[4] ;
    input \SLO_buf[14] ;
    output \spi_data_out_r_39__N_5105[0] ;
    input \SLO_buf[3] ;
    input \SLO_buf[9] ;
    output \spi_data_out_r_39__N_5105[35] ;
    input \SLO_buf[2] ;
    input \SLO_buf[8] ;
    output \spi_data_out_r_39__N_5105[34] ;
    input \SLO_buf[1] ;
    input \SLO_buf[7] ;
    output \spi_data_out_r_39__N_5105[33] ;
    input [31:0]quad_buffer_adj_650;
    input [31:0]quad_count_adj_651;
    output \spi_data_out_r_39__N_1553[0] ;
    output \spi_data_out_r_39__N_1553[31] ;
    input \SLO_buf[0] ;
    input \SLO_buf[6] ;
    output \spi_data_out_r_39__N_5105[32] ;
    input \SLO_buf[19] ;
    input \SLO_buf[29] ;
    output \spi_data_out_r_39__N_5105[15] ;
    output \spi_data_out_r_39__N_1553[30] ;
    output \spi_data_out_r_39__N_1553[29] ;
    output \spi_data_out_r_39__N_1553[28] ;
    output \spi_data_out_r_39__N_1553[27] ;
    input \SLO_buf[18] ;
    input \SLO_buf[28] ;
    output \spi_data_out_r_39__N_5105[14] ;
    output \spi_data_out_r_39__N_1553[26] ;
    input \SLO_buf[17] ;
    input \SLO_buf[27] ;
    output \spi_data_out_r_39__N_5105[13] ;
    output \spi_data_out_r_39__N_2023[25] ;
    output \spi_data_out_r_39__N_1553[25] ;
    output \spi_data_out_r_39__N_1553[24] ;
    input \SLO_buf[16] ;
    input \SLO_buf[26] ;
    output \spi_data_out_r_39__N_5105[12] ;
    output \spi_data_out_r_39__N_1553[23] ;
    input \SLO_buf[15] ;
    input \SLO_buf[25] ;
    output \spi_data_out_r_39__N_5105[11] ;
    input \SLO_buf[24] ;
    output \spi_data_out_r_39__N_5105[10] ;
    output \spi_data_out_r_39__N_1553[22] ;
    input \SLO_buf[13] ;
    input \SLO_buf[23] ;
    output \spi_data_out_r_39__N_5105[9] ;
    output \spi_data_out_r_39__N_1553[21] ;
    output \spi_data_out_r_39__N_1553[20] ;
    output \spi_data_out_r_39__N_1553[19] ;
    output \spi_data_out_r_39__N_1553[18] ;
    output \spi_data_out_r_39__N_1553[17] ;
    output \spi_data_out_r_39__N_1553[16] ;
    output \spi_data_out_r_39__N_1083[16] ;
    output \spi_data_out_r_39__N_1553[15] ;
    output \spi_data_out_r_39__N_1553[14] ;
    output \spi_data_out_r_39__N_1553[13] ;
    output \spi_data_out_r_39__N_1083[15] ;
    input \SLO_buf[12] ;
    input \SLO_buf[22] ;
    output \spi_data_out_r_39__N_5105[8] ;
    output \spi_data_out_r_39__N_1553[12] ;
    input \SLO_buf[11] ;
    input \SLO_buf[21] ;
    output \spi_data_out_r_39__N_5105[7] ;
    output \spi_data_out_r_39__N_1553[11] ;
    input \SLO_buf[10] ;
    input \SLO_buf[20] ;
    output \spi_data_out_r_39__N_5105[6] ;
    output \spi_data_out_r_39__N_5105[5] ;
    output \spi_data_out_r_39__N_1553[10] ;
    output \spi_data_out_r_39__N_5105[4] ;
    output \spi_data_out_r_39__N_1553[9] ;
    output \spi_data_out_r_39__N_1553[8] ;
    output \spi_data_out_r_39__N_1553[7] ;
    output \spi_data_out_r_39__N_1553[6] ;
    output \spi_data_out_r_39__N_5105[3] ;
    output \spi_data_out_r_39__N_1553[5] ;
    output \spi_data_out_r_39__N_1553[4] ;
    output \spi_data_out_r_39__N_1553[3] ;
    output \spi_data_out_r_39__N_2023[18] ;
    output \spi_data_out_r_39__N_1553[2] ;
    output \spi_data_out_r_39__N_1553[1] ;
    output n47_adj_596;
    output \spi_data_out_r_39__N_5105[2] ;
    input \SLO_buf[5] ;
    output \spi_data_out_r_39__N_5105[1] ;
    output spi_data_out_r_39__N_2338;
    output n47_adj_597;
    output \spi_data_out_r_39__N_1083[14] ;
    output \spi_data_out_r_39__N_1083[13] ;
    output n30102;
    input \SLO_buf[4]_adj_598 ;
    input \SLO_buf[14]_adj_599 ;
    output \spi_data_out_r_39__N_4419[0] ;
    input \SLO_buf[3]_adj_600 ;
    input \SLO_buf[9]_adj_601 ;
    output \spi_data_out_r_39__N_4419[35] ;
    output spi_data_out_r_39__N_4505;
    output \spi_data_out_r_39__N_2023[17] ;
    output \spi_data_out_r_39__N_2023[16] ;
    output \spi_data_out_r_39__N_1083[7] ;
    output \spi_data_out_r_39__N_1083[6] ;
    output \spi_data_out_r_39__N_1083[20] ;
    output \spi_data_out_r_39__N_2023[15] ;
    input \status_cntr[12] ;
    output n25212;
    input \SLO_buf[2]_adj_602 ;
    input \SLO_buf[8]_adj_603 ;
    output \spi_data_out_r_39__N_4419[34] ;
    output \spi_data_out_r_39__N_2023[14] ;
    input \SLO_buf[1]_adj_604 ;
    input \SLO_buf[7]_adj_605 ;
    output \spi_data_out_r_39__N_4419[33] ;
    input \SLO_buf[0]_adj_606 ;
    input \SLO_buf[6]_adj_607 ;
    output \spi_data_out_r_39__N_4419[32] ;
    output clear_intrpt_N_3072;
    output \spi_data_out_r_39__N_2023[13] ;
    input \SLO_buf[19]_adj_608 ;
    input \SLO_buf[29]_adj_609 ;
    output \spi_data_out_r_39__N_4419[15] ;
    output \spi_data_out_r_39__N_1083[5] ;
    output \spi_data_out_r_39__N_1083[4] ;
    output \spi_data_out_r_39__N_2023[12] ;
    input \SLO_buf[18]_adj_610 ;
    input \SLO_buf[28]_adj_611 ;
    output \spi_data_out_r_39__N_4419[14] ;
    input \SLO_buf[17]_adj_612 ;
    input \SLO_buf[27]_adj_613 ;
    output \spi_data_out_r_39__N_4419[13] ;
    output \spi_data_out_r_39__N_1083[12] ;
    output spi_data_out_r_39__N_4848;
    output \spi_data_out_r_39__N_1083[3] ;
    output \spi_data_out_r_39__N_1083[2] ;
    output \spi_data_out_r_39__N_2023[11] ;
    input \SLO_buf[16]_adj_614 ;
    input \SLO_buf[26]_adj_615 ;
    output \spi_data_out_r_39__N_4419[12] ;
    output \spi_data_out_r_39__N_2023[10] ;
    input \SLO_buf[15]_adj_616 ;
    input \SLO_buf[25]_adj_617 ;
    output \spi_data_out_r_39__N_4419[11] ;
    input \SLO_buf[24]_adj_618 ;
    output \spi_data_out_r_39__N_4419[10] ;
    input \SLO_buf[13]_adj_619 ;
    input \SLO_buf[23]_adj_620 ;
    output \spi_data_out_r_39__N_4419[9] ;
    input \SLO_buf[12]_adj_621 ;
    input \SLO_buf[22]_adj_622 ;
    output \spi_data_out_r_39__N_4419[8] ;
    input n25885;
    input n30087;
    input \quad_homing[1] ;
    output n1;
    output clk_enable_686;
    output clk_enable_260;
    input clear_intrpt_adj_623;
    output intrpt_out_N_2642;
    output intrpt_out_N_3068;
    output clk_enable_263;
    output clk_enable_807;
    input n12467;
    input n20647;
    input n18654;
    output n12435;
    input n26873;
    output clk_enable_320;
    input n25877;
    input n30075;
    input \quad_homing[1]_adj_624 ;
    output n1_adj_625;
    input n30199;
    input n26821;
    output clk_enable_684;
    input n26089;
    input n26091;
    output clk_enable_255;
    input EM_STOP;
    output clk_enable_23;
    input n26947;
    output clk_enable_253;
    input pwm_out_N_3169;
    input pwm_out_N_3153;
    output clk_enable_15;
    input n26107;
    output n26113;
    input clear_intrpt_adj_626;
    output intrpt_out_N_2997;
    output clk_enable_687;
    input n30045;
    output clk_enable_759;
    output clk_enable_727;
    input n11008;
    input pwm_out_1_N_6491;
    output clk_enable_613;
    input n26957;
    output clk_enable_520;
    output clk_enable_232;
    output clk_enable_28;
    output clk_enable_226;
    output clk_enable_639;
    input pwm_out_3_N_6530;
    output clk_enable_1105;
    input pwm_out_4_N_6549;
    output clk_enable_1107;
    output clk_enable_757;
    output clk_enable_245;
    input pwm_out_2_N_6511;
    output clk_enable_22;
    output clk_enable_488;
    input n26633;
    output clk_enable_641;
    output clk_enable_638;
    output clk_enable_959;
    output clk_enable_235;
    output intrpt_out_N_2713;
    output n57;
    input reset_r_N_4129;
    output clk_enable_761;
    output n29998;
    output clk_enable_738;
    input n25881;
    input n30095;
    input \quad_homing[1]_adj_627 ;
    output n1_adj_628;
    output clk_enable_652;
    input quad_set_valid_N_2098;
    output clk_enable_683;
    output clk_enable_211;
    output n2109;
    input n25893;
    input n30055;
    input \quad_homing[1]_adj_629 ;
    output n1_adj_630;
    input n25869;
    input n30043;
    input \quad_homing[1]_adj_631 ;
    output n1_adj_632;
    input n25873;
    input n30091;
    input \quad_homing[1]_adj_633 ;
    output n1_adj_634;
    input n28476;
    output clk_enable_32;
    output intrpt_out_N_2855;
    output clk_enable_178;
    output intrpt_out_N_2784;
    output clk_enable_842;
    output clk_enable_627;
    output clk_enable_234;
    input quad_set_valid_N_2333;
    output clk_enable_315;
    input \SLO_buf[11]_adj_635 ;
    input \SLO_buf[21]_adj_636 ;
    output \spi_data_out_r_39__N_4419[7] ;
    input clk_enable_256;
    input n29999;
    output clk_enable_12;
    output clk_enable_749;
    output clk_enable_388;
    input n26207;
    output clk_enable_898;
    output clk_enable_180;
    input n18_adj_637;
    output n2193;
    input \SLO_buf[10]_adj_638 ;
    input \SLO_buf[20]_adj_639 ;
    output \spi_data_out_r_39__N_4419[6] ;
    output clk_enable_244;
    output intrpt_out_N_2926;
    input pwm_out_1_N_6306;
    output clk_100k_enable_1;
    input n25889;
    input n30083;
    input \quad_homing[1]_adj_640 ;
    output n1_adj_641;
    output clk_enable_595;
    output n30039;
    output \spi_data_out_r_39__N_2023[9] ;
    output \spi_data_out_r_39__N_1083[24] ;
    output clear_intrpt_N_3001;
    output \spi_data_out_r_39__N_2023[8] ;
    output \spi_data_out_r_39__N_1083[11] ;
    output \spi_data_out_r_39__N_2023[7] ;
    output \spi_data_out_r_39__N_1083[27] ;
    output \spi_data_out_r_39__N_4419[5] ;
    output \spi_data_out_r_39__N_4419[4] ;
    output \spi_data_out_r_39__N_2023[6] ;
    output n27095;
    output spi_data_out_r_39__N_1868;
    output n29992;
    output \spi_data_out_r_39__N_4419[3] ;
    output \spi_data_out_r_39__N_2023[5] ;
    output \spi_data_out_r_39__N_2023[24] ;
    output \spi_data_out_r_39__N_4419[2] ;
    output spi_data_out_r_39__N_5191;
    output spi_data_out_r_39__N_5534;
    output spi_data_out_r_39__N_5877;
    output \spi_data_out_r_39__N_1083[23] ;
    output spi_data_out_r_39__N_6220;
    output \spi_data_out_r_39__N_2023[4] ;
    output \spi_data_out_r_39__N_2023[23] ;
    output \spi_data_out_r_39__N_1083[1] ;
    output \spi_data_out_r_39__N_1083[26] ;
    output spi_data_out_r_39__N_1398;
    output \spi_data_out_r_39__N_1083[25] ;
    output \spi_data_out_r_39__N_1083[30] ;
    output n30013;
    output \spi_data_out_r_39__N_2023[3] ;
    input \SLO_buf[5]_adj_642 ;
    output \spi_data_out_r_39__N_4419[1] ;
    output \spi_data_out_r_39__N_2023[2] ;
    output \spi_data_out_r_39__N_2023[1] ;
    output \spi_data_out_r_39__N_1083[10] ;
    output \spi_data_out_r_39__N_2023[0] ;
    output \spi_data_out_r_39__N_2023[22] ;
    input n30007;
    output clk_enable_38;
    output \spi_data_out_r_39__N_2023[21] ;
    output n30020;
    output \spi_data_out_r_39__N_2023[31] ;
    output clk_enable_227;
    output \spi_data_out_r_39__N_2023[30] ;
    output \spi_data_out_r_39__N_2023[29] ;
    output \spi_data_out_r_39__N_1083[28] ;
    output \spi_data_out_r_39__N_2023[28] ;
    output \spi_data_out_r_39__N_2023[27] ;
    output \spi_data_out_r_39__N_1083[21] ;
    input n22554;
    input pwm;
    input n4_adj_643;
    input \status_cntr[11] ;
    output \spi_data_out_r_39__N_1083[0] ;
    output spi_data_out_r_39__N_2103;
    output spi_data_out_r_39__N_1163;
    output \spi_data_out_r_39__N_2493[0] ;
    output \spi_data_out_r_39__N_2493[31] ;
    output \spi_data_out_r_39__N_2493[30] ;
    output spi_data_out_r_39__N_1633;
    output spi_data_out_r_39__N_2573;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire spi_clk_i /* synthesis is_clock=1 */ ;   // c:/s_links/sources/config_hex/ip/spi_slave_efb.v(34[10:19])
    
    wire clk_enable_624;
    wire [7:0]spi_addr;   // c:/s_links/sources/mcm_top.v(80[28:36])
    
    wire spi_sdo_valid, spi_sdo_valid_N_296, clk_enable_48;
    wire [39:0]spi_data;   // c:/s_links/sources/spi_slave_top.v(70[23:31])
    
    wire spi_scsn_dly, n30142, clk_enable_776;
    wire [15:0]spi_cmd;   // c:/s_links/sources/mcm_top.v(79[27:34])
    wire [39:0]spi_sdo;   // c:/s_links/sources/spi_slave_top.v(74[23:30])
    
    wire n8400, clk_enable_228, spi_addr_valid_r_N_303, n28396, n26563;
    wire [39:0]spi_sdo_r;   // c:/s_links/sources/spi_slave_top.v(66[23:32])
    
    wire clk_enable_963, n23424, n30022, n30033, n28514, n28398, 
        n25833, n24065, n28494, n28540;
    wire [39:0]mem_rdata_7__N_185;
    
    wire n26515, n33, n28516, n26921, n20598, n26923, n26919;
    wire [39:0]spi_sdo_39__N_145;
    
    wire n26911, n26917, n26907, n26905, n26895, n26897, n26893, 
        n26885, n26891, n26881, n26879, n26755, n26757, n26753, 
        n26727, n26745, n26729, n26723, n26749, n26737, n26739, 
        n26733, n30016, n28526, n28488, n25983, n25993, n28518, 
        n30141, n30140, n26539, n26047, n26059, n26587, n30150, 
        n26843, n28448, n26841, n26701, n25380, n28298, n26689, 
        n28452, n28304, n28450, n26667, n28492, n25671, n26063, 
        n28498, n26033, n28364, n28336, n26219, n26233, n30139, 
        n26249, n28366, n26023, n25853, n26075, n26077;
    wire [7:0]mem_rdata;   // c:/s_links/sources/spi_slave_top.v(64[32:41])
    
    wire n23427, n23429, n23425, n30010, n26415, clk_enable_961, 
        n23426, n23430, n23423, n23428, n30011, n30036, wb_cyc_i, 
        clk_enable_172;
    wire [7:0]wb_adr_i;   // c:/s_links/sources/spi_slave_top.v(47[44:52])
    wire [7:0]address;   // c:/s_links/sources/spi_slave_top.v(52[44:51])
    
    wire wb_we_i, wb_we_i_N_344;
    wire [7:0]wb_dat_i;   // c:/s_links/sources/spi_slave_top.v(48[44:52])
    wire [7:0]wr_data;   // c:/s_links/sources/spi_slave_top.v(54[44:51])
    
    wire wb_sm, spi_cmd_start;
    wire [7:0]address_7__N_549;
    wire [7:0]address_7__N_565;
    
    wire wr_en, wr_en_N_355, rd_en, n29;
    wire [7:0]wb_dat_o;   // c:/s_links/sources/spi_slave_top.v(49[44:52])
    
    FD1P3IX spi_addr_r__i0 (.D(spi_addr[0]), .SP(clk_enable_624), .CD(n30080), 
            .CK(clk), .Q(spi_addr_r[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i0.GSR = "DISABLED";
    FD1S3IX spi_sdo_valid_52 (.D(spi_sdo_valid_N_296), .CK(clk), .CD(n30185), 
            .Q(spi_sdo_valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo_valid_52.GSR = "DISABLED";
    FD1P3IX spi_data_valid_r_58 (.D(spi_data_valid), .SP(clk_enable_48), 
            .CD(n30080), .CK(clk), .Q(spi_data_valid_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_valid_r_58.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_635 (.A(n23916), .B(spi_addr_r[3]), .Z(n30035)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_635.init = 16'h2222;
    FD1P3IX spi_data_r__i0 (.D(spi_data[0]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i0.GSR = "DISABLED";
    FD1S3IX spi_scsn_dly_59 (.D(spi_scsn_c), .CK(clk), .CD(n30185), .Q(spi_scsn_dly)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(153[9] 158[5])
    defparam spi_scsn_dly_59.GSR = "DISABLED";
    LUT4 i24023_2_lut (.A(spi_addr_valid), .B(spi_cmd_valid), .Z(clk_enable_48)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/spi_slave_top.v(137[8] 149[6])
    defparam i24023_2_lut.init = 16'hdddd;
    FD1P3IX spi_data_r__i31 (.D(spi_data[31]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i31.GSR = "DISABLED";
    FD1P3IX spi_data_r__i30 (.D(spi_data[30]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i30.GSR = "DISABLED";
    FD1P3IX spi_data_r__i29 (.D(spi_data[29]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i29.GSR = "DISABLED";
    FD1P3IX spi_data_r__i28 (.D(spi_data[28]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i28.GSR = "DISABLED";
    FD1P3IX spi_data_r__i27 (.D(spi_data[27]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i27.GSR = "DISABLED";
    FD1P3IX spi_data_r__i26 (.D(spi_data[26]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i26.GSR = "DISABLED";
    FD1P3IX spi_data_r__i25 (.D(spi_data[25]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i25.GSR = "DISABLED";
    FD1P3IX spi_data_r__i24 (.D(spi_data[24]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i24.GSR = "DISABLED";
    FD1P3IX spi_data_r__i23 (.D(spi_data[23]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i23.GSR = "DISABLED";
    FD1P3IX spi_data_r__i22 (.D(spi_data[22]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i22.GSR = "DISABLED";
    FD1P3IX spi_data_r__i21 (.D(spi_data[21]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i21.GSR = "DISABLED";
    FD1P3IX spi_data_r__i20 (.D(spi_data[20]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i20.GSR = "DISABLED";
    FD1P3IX spi_data_r__i19 (.D(spi_data[19]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i19.GSR = "DISABLED";
    FD1P3IX spi_data_r__i18 (.D(spi_data[18]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i18.GSR = "DISABLED";
    FD1P3IX spi_data_r__i17 (.D(spi_data[17]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i17.GSR = "DISABLED";
    FD1P3IX spi_data_r__i16 (.D(spi_data[16]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i16.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(n30142), .B(spi_cmd_r[1]), .C(n28328), .D(spi_addr_r[0]), 
         .Z(n26327)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_3_lut_4_lut.init = 16'h0008;
    FD1P3IX spi_data_r__i15 (.D(spi_data[15]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i15.GSR = "DISABLED";
    FD1P3IX spi_data_r__i14 (.D(spi_data[14]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i14.GSR = "DISABLED";
    FD1P3IX spi_data_r__i13 (.D(spi_data[13]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i13.GSR = "DISABLED";
    FD1P3IX spi_data_r__i12 (.D(spi_data[12]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i12.GSR = "DISABLED";
    FD1P3IX spi_data_r__i11 (.D(spi_data[11]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i11.GSR = "DISABLED";
    FD1P3IX spi_data_r__i10 (.D(spi_data[10]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i10.GSR = "DISABLED";
    FD1P3IX spi_data_r__i9 (.D(spi_data[9]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i9.GSR = "DISABLED";
    FD1P3IX spi_data_r__i8 (.D(spi_data[8]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i8.GSR = "DISABLED";
    FD1P3IX spi_data_r__i7 (.D(spi_data[7]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i7.GSR = "DISABLED";
    FD1P3IX spi_data_r__i6 (.D(spi_data[6]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i6.GSR = "DISABLED";
    FD1P3IX spi_data_r__i5 (.D(spi_data[5]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i5.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i0 (.D(spi_cmd[0]), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i0.GSR = "DISABLED";
    FD1P3IX spi_data_r__i4 (.D(spi_data[4]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i4.GSR = "DISABLED";
    FD1P3IX spi_data_r__i3 (.D(spi_data[3]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i3.GSR = "DISABLED";
    FD1P3IX spi_data_r__i2 (.D(spi_data[2]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i2.GSR = "DISABLED";
    FD1P3IX spi_data_r__i1 (.D(spi_data[1]), .SP(clk_enable_161), .CD(n30080), 
            .CK(clk), .Q(\spi_data_r[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i1.GSR = "DISABLED";
    FD1P3IX spi_sdo__i0 (.D(\spi_data_out_r[0] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i0.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_744 (.A(n30142), .B(spi_cmd_r[1]), .C(n26621), 
         .D(spi_addr_r[0]), .Z(n26819)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_3_lut_4_lut_adj_744.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n30142), .B(spi_cmd_r[1]), .C(n27013), 
         .D(spi_cmd_r[3]), .Z(n27015)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i23822_3_lut_4_lut (.A(n30144), .B(spi_addr_r[2]), .C(n30155), 
         .D(n18440), .Z(n28524)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23822_3_lut_4_lut.init = 16'hfffe;
    FD1P3IX spi_addr_valid_r_56 (.D(spi_addr_valid_r_N_303), .SP(clk_enable_228), 
            .CD(n30080), .CK(clk), .Q(spi_sdo_valid_N_296)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_valid_r_56.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(spi_cmd_r[2]), .B(n4), .C(spi_cmd_r[3]), .D(n30044), 
         .Z(n23526)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_4_lut.init = 16'h0400;
    LUT4 i1_4_lut_adj_745 (.A(n30044), .B(n26545), .C(n28396), .D(spi_addr_r[3]), 
         .Z(n26563)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_745.init = 16'h0008;
    LUT4 i23694_2_lut (.A(spi_cmd_r[3]), .B(spi_addr_r[1]), .Z(n28396)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23694_2_lut.init = 16'heeee;
    FD1P3AX spi_sdo_r__i0 (.D(n23424), .SP(clk_enable_963), .CK(clk), 
            .Q(spi_sdo_r[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i0.GSR = "DISABLED";
    LUT4 i23828_2_lut_rep_622_4_lut (.A(n30155), .B(n30144), .C(spi_addr_r[2]), 
         .D(spi_addr_r[0]), .Z(n30022)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23828_2_lut_rep_622_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_633_4_lut (.A(n30155), .B(n30144), .C(spi_addr_r[2]), 
         .D(spi_addr_r[0]), .Z(n30033)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_633_4_lut.init = 16'h0100;
    LUT4 i23812_2_lut_3_lut_4_lut (.A(spi_addr_r[0]), .B(n30155), .C(spi_addr_r[2]), 
         .D(n30144), .Z(n28514)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23812_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_746 (.A(n28398), .B(n30151), .C(n30094), .D(spi_addr_r[0]), 
         .Z(n25833)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_746.init = 16'h0004;
    LUT4 i1_4_lut_adj_747 (.A(spi_cmd_r[0]), .B(n24065), .C(spi_cmd_r[2]), 
         .D(n30044), .Z(quad_set_valid_N_1158)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_4_lut_adj_747.init = 16'h0400;
    LUT4 i1_4_lut_adj_748 (.A(n28494), .B(n23916), .C(n28396), .D(spi_addr_r[0]), 
         .Z(n24065)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_748.init = 16'h0004;
    FD1P3IX spi_addr_r__i7 (.D(spi_addr[7]), .SP(clk_enable_624), .CD(n30080), 
            .CK(clk), .Q(spi_addr_r[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i7.GSR = "DISABLED";
    FD1P3IX spi_addr_r__i6 (.D(spi_addr[6]), .SP(clk_enable_624), .CD(n30080), 
            .CK(clk), .Q(spi_addr_r[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i6.GSR = "DISABLED";
    FD1P3IX spi_addr_r__i5 (.D(spi_addr[5]), .SP(clk_enable_624), .CD(n30080), 
            .CK(clk), .Q(spi_addr_r[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i5.GSR = "DISABLED";
    FD1P3IX spi_addr_r__i4 (.D(spi_addr[4]), .SP(clk_enable_624), .CD(n30080), 
            .CK(clk), .Q(spi_addr_r[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i4.GSR = "DISABLED";
    FD1P3IX spi_addr_r__i3 (.D(spi_addr[3]), .SP(clk_enable_624), .CD(n30080), 
            .CK(clk), .Q(spi_addr_r[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i3.GSR = "DISABLED";
    FD1P3IX spi_addr_r__i2 (.D(spi_addr[2]), .SP(clk_enable_624), .CD(n30080), 
            .CK(clk), .Q(spi_addr_r[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i2.GSR = "DISABLED";
    FD1P3IX spi_addr_r__i1 (.D(spi_addr[1]), .SP(clk_enable_624), .CD(n30080), 
            .CK(clk), .Q(spi_addr_r[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i1.GSR = "DISABLED";
    LUT4 i23838_4_lut (.A(n30094), .B(n23732), .C(n28398), .D(spi_addr_r[0]), 
         .Z(n28540)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23838_4_lut.init = 16'hfffe;
    LUT4 mux_18_i32_3_lut (.A(spi_sdo_r[23]), .B(spi_sdo[31]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i32_3_lut.init = 16'hcaca;
    LUT4 mux_18_i36_3_lut (.A(spi_sdo_r[27]), .B(spi_sdo[35]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[35])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i36_3_lut.init = 16'hcaca;
    LUT4 mux_18_i39_3_lut (.A(spi_sdo_r[30]), .B(spi_sdo[38]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[38])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i39_3_lut.init = 16'hcaca;
    LUT4 mux_18_i33_3_lut (.A(spi_sdo_r[24]), .B(spi_sdo[32]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[32])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i33_3_lut.init = 16'hcaca;
    LUT4 mux_18_i37_3_lut (.A(spi_sdo_r[28]), .B(spi_sdo[36]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[36])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i37_3_lut.init = 16'hcaca;
    LUT4 mux_18_i40_3_lut (.A(spi_sdo_r[31]), .B(spi_sdo[39]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[39])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i40_3_lut.init = 16'hcaca;
    LUT4 mux_18_i30_3_lut (.A(spi_sdo_r[21]), .B(spi_sdo[29]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i30_3_lut.init = 16'hcaca;
    LUT4 mux_18_i34_3_lut (.A(spi_sdo_r[25]), .B(spi_sdo[33]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[33])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i34_3_lut.init = 16'hcaca;
    LUT4 mux_18_i31_3_lut (.A(spi_sdo_r[22]), .B(spi_sdo[30]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i31_3_lut.init = 16'hcaca;
    LUT4 mux_18_i35_3_lut (.A(spi_sdo_r[26]), .B(spi_sdo[34]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[34])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i35_3_lut.init = 16'hcaca;
    LUT4 mux_18_i38_3_lut (.A(spi_sdo_r[29]), .B(spi_sdo[37]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[37])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i38_3_lut.init = 16'hcaca;
    LUT4 i23696_2_lut (.A(spi_addr_r[2]), .B(spi_addr_r[1]), .Z(n28398)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23696_2_lut.init = 16'heeee;
    LUT4 mux_18_i20_3_lut (.A(spi_sdo_r[11]), .B(spi_sdo[19]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i20_3_lut.init = 16'hcaca;
    LUT4 mux_18_i24_3_lut (.A(spi_sdo_r[15]), .B(spi_sdo[23]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i24_3_lut.init = 16'hcaca;
    LUT4 mux_18_i27_3_lut (.A(spi_sdo_r[18]), .B(spi_sdo[26]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i27_3_lut.init = 16'hcaca;
    LUT4 mux_18_i21_3_lut (.A(spi_sdo_r[12]), .B(spi_sdo[20]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i21_3_lut.init = 16'hcaca;
    LUT4 mux_18_i25_3_lut (.A(spi_sdo_r[16]), .B(spi_sdo[24]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i25_3_lut.init = 16'hcaca;
    LUT4 mux_18_i28_3_lut (.A(spi_sdo_r[19]), .B(spi_sdo[27]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i28_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_749 (.A(n26497), .B(n30044), .C(n30209), .D(spi_addr_r[2]), 
         .Z(n26515)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_749.init = 16'h0008;
    LUT4 i23814_4_lut (.A(n33), .B(n28260), .C(spi_addr_r[0]), .D(n30214), 
         .Z(n28516)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23814_4_lut.init = 16'hfffe;
    LUT4 mux_18_i18_3_lut (.A(spi_sdo_r[9]), .B(spi_sdo[17]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i18_3_lut.init = 16'hcaca;
    FD1P3IX spi_cmd_r__i1 (.D(spi_cmd[1]), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i1.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i2 (.D(\spi_cmd[2] ), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i2.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i3 (.D(spi_cmd[3]), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i3.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i4 (.D(spi_cmd[4]), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i4.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i5 (.D(spi_cmd[5]), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i5.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i6 (.D(spi_cmd[6]), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i6.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i7 (.D(spi_cmd[7]), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i7.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i8 (.D(spi_cmd[8]), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i8.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i9 (.D(spi_cmd[9]), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i9.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i10 (.D(spi_cmd[10]), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i10.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i11 (.D(spi_cmd[11]), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i11.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i12 (.D(spi_cmd[12]), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i12.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i13 (.D(spi_cmd[13]), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i13.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i14 (.D(spi_cmd[14]), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i14.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i15 (.D(spi_cmd[15]), .SP(clk_enable_776), .CD(n30080), 
            .CK(clk), .Q(spi_cmd_r[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i15.GSR = "DISABLED";
    FD1P3IX spi_sdo__i1 (.D(\spi_data_out_r[1] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i1.GSR = "DISABLED";
    LUT4 i51_2_lut (.A(\spi_data_r[16] ), .B(\spi_data_r[17] ), .Z(n33)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i51_2_lut.init = 16'heeee;
    LUT4 mux_18_i22_3_lut (.A(spi_sdo_r[13]), .B(spi_sdo[21]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i22_3_lut.init = 16'hcaca;
    LUT4 mux_18_i19_3_lut (.A(spi_sdo_r[10]), .B(spi_sdo[18]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i19_3_lut.init = 16'hcaca;
    LUT4 mux_18_i23_3_lut (.A(spi_sdo_r[14]), .B(spi_sdo[22]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i23_3_lut.init = 16'hcaca;
    LUT4 mux_18_i26_3_lut (.A(spi_sdo_r[17]), .B(spi_sdo[25]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i26_3_lut.init = 16'hcaca;
    LUT4 mux_18_i29_3_lut (.A(spi_sdo_r[20]), .B(spi_sdo[28]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i29_3_lut.init = 16'hcaca;
    LUT4 mux_18_i12_3_lut (.A(spi_sdo_r[3]), .B(spi_sdo[11]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i12_3_lut.init = 16'hcaca;
    LUT4 mux_18_i15_3_lut (.A(spi_sdo_r[6]), .B(spi_sdo[14]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i15_3_lut.init = 16'hcaca;
    LUT4 mux_18_i9_3_lut (.A(spi_sdo_r[0]), .B(spi_sdo[8]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i9_3_lut.init = 16'hcaca;
    LUT4 mux_18_i13_3_lut (.A(spi_sdo_r[4]), .B(spi_sdo[12]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i13_3_lut.init = 16'hcaca;
    LUT4 mux_18_i16_3_lut (.A(spi_sdo_r[7]), .B(spi_sdo[15]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i16_3_lut.init = 16'hcaca;
    LUT4 mux_18_i10_3_lut (.A(spi_sdo_r[1]), .B(spi_sdo[9]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i10_3_lut.init = 16'hcaca;
    LUT4 mux_18_i11_3_lut (.A(spi_sdo_r[2]), .B(spi_sdo[10]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i11_3_lut.init = 16'hcaca;
    LUT4 mux_18_i14_3_lut (.A(spi_sdo_r[5]), .B(spi_sdo[13]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i14_3_lut.init = 16'hcaca;
    LUT4 mux_18_i17_3_lut (.A(spi_sdo_r[8]), .B(spi_sdo[16]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i17_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_750 (.A(n26921), .B(n20598), .C(n26923), .D(n26919), 
         .Z(spi_sdo_39__N_145[8])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_750.init = 16'hfffe;
    FD1P3IX spi_sdo__i3 (.D(\spi_data_out_r[3] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i3.GSR = "DISABLED";
    FD1P3IX spi_sdo__i4 (.D(\spi_data_out_r[4] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i4.GSR = "DISABLED";
    FD1P3IX spi_sdo__i5 (.D(\spi_data_out_r[5] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i5.GSR = "DISABLED";
    FD1P3IX spi_sdo__i6 (.D(\spi_data_out_r[6] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i6.GSR = "DISABLED";
    FD1P3IX spi_sdo__i7 (.D(\spi_data_out_r[7] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i7.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_751 (.A(\spi_data_out_r_39__N_5197[8] ), .B(n26911), 
         .C(n16), .D(spi_data_out_r_39__N_5237), .Z(n26921)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_751.init = 16'hfefc;
    FD1P3IX spi_sdo__i10 (.D(\spi_data_out_r[10] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i10.GSR = "DISABLED";
    FD1P3IX spi_sdo__i11 (.D(\spi_data_out_r[11] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i11.GSR = "DISABLED";
    FD1P3IX spi_sdo__i12 (.D(\spi_data_out_r[12] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i12.GSR = "DISABLED";
    FD1P3IX spi_sdo__i13 (.D(\spi_data_out_r[13] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i13.GSR = "DISABLED";
    FD1P3IX spi_sdo__i14 (.D(\spi_data_out_r[14] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i14.GSR = "DISABLED";
    FD1P3IX spi_sdo__i15 (.D(\spi_data_out_r[15] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i15.GSR = "DISABLED";
    FD1P3IX spi_sdo__i16 (.D(\spi_data_out_r[16] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i16.GSR = "DISABLED";
    FD1P3IX spi_sdo__i17 (.D(\spi_data_out_r[17] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i17.GSR = "DISABLED";
    FD1P3IX spi_sdo__i18 (.D(\spi_data_out_r[18] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i18.GSR = "DISABLED";
    FD1P3IX spi_sdo__i19 (.D(\spi_data_out_r[19] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i19.GSR = "DISABLED";
    FD1P3IX spi_sdo__i20 (.D(\spi_data_out_r[20] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i20.GSR = "DISABLED";
    FD1P3IX spi_sdo__i21 (.D(\spi_data_out_r[21] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i21.GSR = "DISABLED";
    FD1P3IX spi_sdo__i22 (.D(\spi_data_out_r[22] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i22.GSR = "DISABLED";
    FD1P3IX spi_sdo__i23 (.D(\spi_data_out_r[23] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i23.GSR = "DISABLED";
    FD1P3IX spi_sdo__i24 (.D(\spi_data_out_r[24] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i24.GSR = "DISABLED";
    FD1P3IX spi_sdo__i25 (.D(\spi_data_out_r[25] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i25.GSR = "DISABLED";
    FD1P3IX spi_sdo__i26 (.D(\spi_data_out_r[26] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i26.GSR = "DISABLED";
    FD1P3IX spi_sdo__i27 (.D(\spi_data_out_r[27] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i27.GSR = "DISABLED";
    FD1P3IX spi_sdo__i28 (.D(\spi_data_out_r[28] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i28.GSR = "DISABLED";
    FD1P3IX spi_sdo__i29 (.D(\spi_data_out_r[29] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i29.GSR = "DISABLED";
    FD1P3IX spi_sdo__i30 (.D(\spi_data_out_r[30] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i30.GSR = "DISABLED";
    FD1P3IX spi_sdo__i31 (.D(\spi_data_out_r[31] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i31.GSR = "DISABLED";
    FD1P3IX spi_sdo__i32 (.D(\spi_data_out_r[32] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i32.GSR = "DISABLED";
    FD1P3IX spi_sdo__i33 (.D(\spi_data_out_r[33] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i33.GSR = "DISABLED";
    FD1P3IX spi_sdo__i34 (.D(\spi_data_out_r[34] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i34.GSR = "DISABLED";
    FD1P3IX spi_sdo__i35 (.D(\spi_data_out_r[35] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i35.GSR = "DISABLED";
    FD1P3IX spi_sdo__i36 (.D(\spi_data_out_r[36] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i36.GSR = "DISABLED";
    FD1P3IX spi_sdo__i37 (.D(\spi_data_out_r[37] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i37.GSR = "DISABLED";
    FD1P3IX spi_sdo__i38 (.D(\spi_data_out_r[38] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i38.GSR = "DISABLED";
    FD1P3IX spi_sdo__i39 (.D(\spi_data_out_r[39] ), .SP(spi_sdo_valid_N_296), 
            .CD(n8400), .CK(clk), .Q(spi_sdo[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i39.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_752 (.A(n26917), .B(\spi_data_out_r_39__N_5540[8] ), 
         .C(n18), .D(spi_data_out_r_39__N_5580), .Z(n26923)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_752.init = 16'hfefa;
    LUT4 i1_4_lut_adj_753 (.A(\spi_data_out_r_39__N_4168[8] ), .B(n26907), 
         .C(n3), .D(spi_data_out_r_39__N_4208), .Z(n26919)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_753.init = 16'hfefc;
    LUT4 i1_4_lut_adj_754 (.A(\spi_data_out_r_39__N_5883[8] ), .B(\spi_data_out_r_39__N_4854[8] ), 
         .C(spi_data_out_r_39__N_5923), .D(spi_data_out_r_39__N_4894), .Z(n26911)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_754.init = 16'heca0;
    LUT4 i1_4_lut_adj_755 (.A(\spi_data_out_r_39__N_2109[8] ), .B(n26905), 
         .C(n5), .D(spi_data_out_r_39__N_2149), .Z(n26917)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_755.init = 16'hfefc;
    LUT4 i1_4_lut_adj_756 (.A(\spi_data_out_r_39__N_1404[8] ), .B(\spi_data_out_r_39__N_934[8] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_974), .Z(n26905)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_756.init = 16'heca0;
    LUT4 i23682_2_lut (.A(spi_addr_r[4]), .B(spi_addr_r[5]), .Z(n28384)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23682_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_757 (.A(\spi_data_out_r_39__N_2344[8] ), .B(\spi_data_out_r_39__N_1874[8] ), 
         .C(spi_data_out_r_39__N_2384), .D(spi_data_out_r_39__N_1914), .Z(n26907)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_757.init = 16'heca0;
    LUT4 i1_4_lut_adj_758 (.A(n26895), .B(n20598), .C(n26897), .D(n26893), 
         .Z(spi_sdo_39__N_145[9])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_758.init = 16'hfffe;
    LUT4 i1_4_lut_adj_759 (.A(\spi_data_out_r_39__N_4168[9] ), .B(n26885), 
         .C(n16_adj_329), .D(spi_data_out_r_39__N_4208), .Z(n26895)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_759.init = 16'hfefc;
    LUT4 i1_4_lut_adj_760 (.A(n26891), .B(\spi_data_out_r_39__N_5883[9] ), 
         .C(n21), .D(spi_data_out_r_39__N_5923), .Z(n26897)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_760.init = 16'hfefa;
    LUT4 i1_4_lut_adj_761 (.A(\spi_data_out_r_39__N_4854[9] ), .B(n26881), 
         .C(n2), .D(spi_data_out_r_39__N_4894), .Z(n26893)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_761.init = 16'hfefc;
    LUT4 i1_4_lut_adj_762 (.A(\spi_data_out_r_39__N_5197[9] ), .B(\spi_data_out_r_39__N_4511[9] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4551), .Z(n26885)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_762.init = 16'heca0;
    LUT4 i1_4_lut_adj_763 (.A(\spi_data_out_r_39__N_1874[9] ), .B(n26879), 
         .C(n5_adj_330), .D(spi_data_out_r_39__N_1914), .Z(n26891)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_763.init = 16'hfefc;
    LUT4 i1_4_lut_adj_764 (.A(\spi_data_out_r_39__N_2344[9] ), .B(\spi_data_out_r_39__N_2109[9] ), 
         .C(spi_data_out_r_39__N_2384), .D(spi_data_out_r_39__N_2149), .Z(n26879)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_764.init = 16'heca0;
    LUT4 i1_4_lut_adj_765 (.A(\spi_data_out_r_39__N_1404[9] ), .B(\spi_data_out_r_39__N_1169[9] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1209), .Z(n26881)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_765.init = 16'heca0;
    LUT4 i1_4_lut_adj_766 (.A(n26755), .B(n20598), .C(n26757), .D(n26753), 
         .Z(spi_sdo_39__N_145[2])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_766.init = 16'hfffe;
    LUT4 i1_4_lut_adj_767 (.A(n26727), .B(n26745), .C(n26729), .D(n26723), 
         .Z(n26755)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_767.init = 16'hfffe;
    LUT4 i1_4_lut_adj_768 (.A(n21_adj_331), .B(n26749), .C(n26737), .D(n19), 
         .Z(n26757)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_768.init = 16'hfffe;
    LUT4 i1_4_lut_adj_769 (.A(\spi_data_out_r_39__N_5197[2] ), .B(n26739), 
         .C(n22), .D(spi_data_out_r_39__N_5237), .Z(n26753)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_769.init = 16'hfefc;
    LUT4 i1_4_lut_adj_770 (.A(\spi_data_out_r_39__N_2863[2] ), .B(\spi_data_out_r_39__N_2721[2] ), 
         .C(clear_intrpt), .D(clear_intrpt_adj_332), .Z(n26727)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_770.init = 16'heca0;
    LUT4 i1_4_lut_adj_771 (.A(\spi_data_out_r_39__N_4511[2] ), .B(\spi_data_out_r_39__N_4168[2] ), 
         .C(spi_data_out_r_39__N_4551), .D(spi_data_out_r_39__N_4208), .Z(n26745)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_771.init = 16'heca0;
    LUT4 i1_4_lut_adj_772 (.A(\spi_data_out_r_39__N_3005[2] ), .B(n14), 
         .C(n9), .D(clear_intrpt_adj_333), .Z(n26729)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_772.init = 16'hfefc;
    LUT4 i1_4_lut_adj_773 (.A(\spi_data_out_r_39__N_2792[2] ), .B(\spi_data_out_r_39__N_2650[2] ), 
         .C(clear_intrpt_adj_334), .D(clear_intrpt_adj_335), .Z(n26723)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_773.init = 16'heca0;
    LUT4 i1_4_lut_adj_774 (.A(\spi_data_out_r_39__N_1169[2] ), .B(n26733), 
         .C(n7), .D(spi_data_out_r_39__N_1209), .Z(n26749)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_774.init = 16'hfefc;
    LUT4 i1_4_lut_adj_775 (.A(\spi_data_out_r_39__N_1639[2] ), .B(\spi_data_out_r_39__N_1404[2] ), 
         .C(spi_data_out_r_39__N_1679), .D(spi_data_out_r_39__N_1444), .Z(n26737)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_775.init = 16'heca0;
    LUT4 i1_4_lut_adj_776 (.A(\spi_data_out_r_39__N_1874[2] ), .B(\spi_data_out_r_39__N_2344[2] ), 
         .C(spi_data_out_r_39__N_1914), .D(spi_data_out_r_39__N_2384), .Z(n26733)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_776.init = 16'heca0;
    LUT4 i1_4_lut_adj_777 (.A(\spi_data_out_r_39__N_3825[2] ), .B(\spi_data_out_r_39__N_934[2] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_974), .Z(n26739)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_777.init = 16'heca0;
    LUT4 i1_4_lut_adj_778 (.A(n30016), .B(n28526), .C(n30151), .D(n28488), 
         .Z(n25721)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_4_lut_adj_778.init = 16'h0020;
    LUT4 i1_4_lut_adj_779 (.A(n25983), .B(n30044), .C(n28358), .D(n30214), 
         .Z(n25993)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_779.init = 16'h0008;
    LUT4 i1_2_lut (.A(spi_addr_r[7]), .B(spi_addr_r[0]), .Z(n25983)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i1_4_lut_adj_780 (.A(n28518), .B(n30151), .C(n30141), .D(n33), 
         .Z(n26435)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_780.init = 16'h0004;
    LUT4 i23816_4_lut (.A(spi_addr_r[0]), .B(n30140), .C(n28384), .D(spi_addr_r[2]), 
         .Z(n28518)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23816_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_781 (.A(n30044), .B(n26521), .C(n28396), .D(spi_addr_r[3]), 
         .Z(n26539)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_781.init = 16'h0008;
    LUT4 i1_4_lut_adj_782 (.A(n30090), .B(spi_cmd_r[4]), .C(spi_addr_r[4]), 
         .D(n26047), .Z(n26059)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_782.init = 16'h0200;
    LUT4 i1_4_lut_adj_783 (.A(n30044), .B(n26569), .C(n28396), .D(spi_addr_r[3]), 
         .Z(n26587)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_783.init = 16'h0008;
    LUT4 i1_4_lut_adj_784 (.A(n30150), .B(n30044), .C(spi_cmd_r[3]), .D(spi_cmd_r[2]), 
         .Z(n26843)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_784.init = 16'h0004;
    LUT4 i1_4_lut_adj_785 (.A(n28448), .B(spi_addr_r[5]), .C(n30140), 
         .D(spi_cmd_r[0]), .Z(n26841)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_785.init = 16'h0100;
    LUT4 i1_4_lut_adj_786 (.A(n26701), .B(n25380), .C(n28448), .D(n28298), 
         .Z(n20598)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_4_lut_adj_786.init = 16'h0008;
    LUT4 i1_4_lut_adj_787 (.A(spi_addr_r[5]), .B(n30140), .C(spi_cmd[15]), 
         .D(spi_addr_r[3]), .Z(n26701)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_787.init = 16'h1000;
    LUT4 i1_4_lut_adj_788 (.A(n26689), .B(n28452), .C(spi_cmd[4]), .D(spi_cmd[9]), 
         .Z(n25380)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_788.init = 16'h0002;
    LUT4 i23596_2_lut (.A(spi_addr_r[2]), .B(\spi_cmd[2] ), .Z(n28298)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23596_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_789 (.A(n28304), .B(spi_cmd[7]), .C(n28450), .D(n26667), 
         .Z(n26689)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_789.init = 16'h0100;
    LUT4 i23602_2_lut (.A(spi_cmd[10]), .B(spi_cmd[5]), .Z(n28304)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23602_2_lut.init = 16'heeee;
    LUT4 i23748_4_lut (.A(spi_cmd[14]), .B(spi_cmd[13]), .C(spi_cmd[12]), 
         .D(spi_cmd[6]), .Z(n28450)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23748_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut (.A(spi_cmd[8]), .B(spi_sdo_valid_N_296), .C(spi_cmd[0]), 
         .Z(n26667)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut.init = 16'h4040;
    LUT4 i1_4_lut_adj_790 (.A(n28492), .B(n24066), .C(n28340), .D(n25671), 
         .Z(quad_set_valid_N_1393)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_790.init = 16'h0400;
    LUT4 i1_4_lut_adj_791 (.A(spi_addr_r[4]), .B(spi_addr_r[2]), .C(n26063), 
         .D(n30142), .Z(n25671)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_791.init = 16'h1000;
    LUT4 i1_2_lut_adj_792 (.A(spi_addr_r[0]), .B(spi_cmd_r[1]), .Z(n26063)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_792.init = 16'h8888;
    LUT4 i1_4_lut_adj_793 (.A(n30016), .B(n28498), .C(n30151), .D(n30071), 
         .Z(n25571)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_4_lut_adj_793.init = 16'h0020;
    LUT4 spi_addr_valid_r_I_5_3_lut (.A(spi_sdo_valid_N_296), .B(spi_addr_valid), 
         .C(spi_data_valid), .Z(spi_addr_valid_r_N_303)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // c:/s_links/sources/mcm_top.v(177[3] 197[2])
    defparam spi_addr_valid_r_I_5_3_lut.init = 16'hecec;
    LUT4 i1_3_lut_adj_794 (.A(spi_cmd_r[4]), .B(spi_cmd_r[2]), .C(spi_cmd_r[1]), 
         .Z(n26033)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut_adj_794.init = 16'h1010;
    LUT4 i23662_2_lut (.A(spi_cmd_r[0]), .B(spi_cmd_r[5]), .Z(n28364)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23662_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_795 (.A(n30155), .B(n28448), .C(n28336), .D(n26219), 
         .Z(n26233)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_795.init = 16'h0100;
    LUT4 i23634_2_lut (.A(spi_addr_r[2]), .B(spi_cmd_r[0]), .Z(n28336)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23634_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_796 (.A(spi_addr_r[6]), .B(spi_cmd_r[2]), .Z(n26219)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_796.init = 16'h4444;
    LUT4 i1_4_lut_adj_797 (.A(n26243), .B(n30139), .C(spi_addr_r[0]), 
         .D(n30155), .Z(n26249)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_797.init = 16'h0002;
    LUT4 i23664_2_lut (.A(spi_cmd_r[0]), .B(spi_cmd_r[4]), .Z(n28366)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23664_2_lut.init = 16'heeee;
    LUT4 i1_3_lut_adj_798 (.A(spi_cmd_r[5]), .B(spi_cmd_r[1]), .C(spi_cmd_r[2]), 
         .Z(n26023)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_3_lut_adj_798.init = 16'h4040;
    LUT4 i1_4_lut_adj_799 (.A(n23916), .B(n30062), .C(spi_addr_r[3]), 
         .D(n25853), .Z(n25859)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_4_lut_adj_799.init = 16'h0800;
    LUT4 i1_2_lut_adj_800 (.A(spi_addr_r[0]), .B(resetn_c), .Z(n25853)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_adj_800.init = 16'h8888;
    LUT4 i23686_2_lut_rep_809 (.A(spi_addr_r[3]), .B(spi_cmd_r[3]), .Z(n30209)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23686_2_lut_rep_809.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(spi_addr_r[3]), .B(spi_cmd_r[3]), .C(n23916), 
         .Z(n24066)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_rep_810 (.A(spi_addr_r[2]), .B(spi_cmd_r[1]), .Z(n30210)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_810.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_801 (.A(spi_addr_r[2]), .B(spi_cmd_r[1]), .C(spi_addr_r[0]), 
         .Z(n26047)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_801.init = 16'h8080;
    LUT4 i23698_2_lut_rep_813 (.A(spi_addr_r[7]), .B(spi_addr_r[4]), .Z(n30213)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23698_2_lut_rep_813.init = 16'heeee;
    LUT4 i1_2_lut_rep_595_4_lut (.A(n23916), .B(n28524), .C(n30023), .D(spi_addr_r[0]), 
         .Z(n29995)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_595_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_rep_596_4_lut (.A(n23916), .B(n28524), .C(n30023), .D(spi_addr_r[0]), 
         .Z(n29996)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_596_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_4_lut (.A(n30016), .B(n23916), .C(n30023), .D(n30033), 
         .Z(clk_enable_254)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_4_lut_adj_802 (.A(n30016), .B(n23916), .C(n30023), .D(n30022), 
         .Z(clk_enable_259)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_4_lut_adj_802.init = 16'h0080;
    LUT4 i1_4_lut_adj_803 (.A(n26075), .B(spi_addr_r[4]), .C(spi_addr_r[2]), 
         .D(spi_cmd_r[4]), .Z(n26077)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_803.init = 16'h0002;
    LUT4 i1_4_lut_adj_804 (.A(spi_cmd_r[5]), .B(n30155), .C(spi_addr_r[6]), 
         .D(n26063), .Z(n26075)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_804.init = 16'h0100;
    FD1P3IX spi_sdo_r__i31 (.D(mem_rdata_7__N_185[31]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i31.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i35 (.D(mem_rdata_7__N_185[35]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(mem_rdata[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i35.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i38 (.D(mem_rdata_7__N_185[38]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(mem_rdata[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i38.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i32 (.D(mem_rdata_7__N_185[32]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(mem_rdata[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i32.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i36 (.D(mem_rdata_7__N_185[36]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(mem_rdata[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i36.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i39 (.D(mem_rdata_7__N_185[39]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(mem_rdata[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i39.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i29 (.D(mem_rdata_7__N_185[29]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i29.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i33 (.D(mem_rdata_7__N_185[33]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(mem_rdata[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i33.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i30 (.D(mem_rdata_7__N_185[30]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i30.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i34 (.D(mem_rdata_7__N_185[34]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(mem_rdata[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i34.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i37 (.D(mem_rdata_7__N_185[37]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(mem_rdata[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i37.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i19 (.D(mem_rdata_7__N_185[19]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i19.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i23 (.D(mem_rdata_7__N_185[23]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i23.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i26 (.D(mem_rdata_7__N_185[26]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i26.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i20 (.D(mem_rdata_7__N_185[20]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i20.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i24 (.D(mem_rdata_7__N_185[24]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i24.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i27 (.D(mem_rdata_7__N_185[27]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i27.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i17 (.D(mem_rdata_7__N_185[17]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i17.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i21 (.D(mem_rdata_7__N_185[21]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i21.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i18 (.D(mem_rdata_7__N_185[18]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i18.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i22 (.D(mem_rdata_7__N_185[22]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i22.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i25 (.D(mem_rdata_7__N_185[25]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i25.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i28 (.D(mem_rdata_7__N_185[28]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i28.GSR = "DISABLED";
    FD1P3AX spi_sdo_r__i7 (.D(n23427), .SP(clk_enable_963), .CK(clk), 
            .Q(spi_sdo_r[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i7.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i11 (.D(mem_rdata_7__N_185[11]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i11.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i14 (.D(mem_rdata_7__N_185[14]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i14.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i8 (.D(mem_rdata_7__N_185[8]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i8.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i12 (.D(mem_rdata_7__N_185[12]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i12.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i15 (.D(mem_rdata_7__N_185[15]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i15.GSR = "DISABLED";
    FD1P3AX spi_sdo_r__i5 (.D(n23429), .SP(clk_enable_963), .CK(clk), 
            .Q(spi_sdo_r[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i5.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i9 (.D(mem_rdata_7__N_185[9]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i9.GSR = "DISABLED";
    FD1P3AX spi_sdo_r__i6 (.D(n23425), .SP(clk_enable_963), .CK(clk), 
            .Q(spi_sdo_r[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i6.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i10 (.D(mem_rdata_7__N_185[10]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i10.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i13 (.D(mem_rdata_7__N_185[13]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i13.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i16 (.D(mem_rdata_7__N_185[16]), .SP(clk_enable_963), 
            .CD(n30185), .CK(clk), .Q(spi_sdo_r[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i16.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_593_3_lut_4_lut (.A(n30070), .B(spi_addr_r[0]), .C(n23526), 
         .D(n30035), .Z(n29993)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_593_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_3_lut_rep_610_4_lut (.A(n30062), .B(spi_addr_r[3]), .C(n28524), 
         .D(n23916), .Z(n30010)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_3_lut_rep_610_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_805 (.A(n30062), .B(spi_addr_r[3]), .C(spi_cmd_r[3]), 
         .D(n30044), .Z(n26415)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_3_lut_4_lut_adj_805.init = 16'h0200;
    FD1P3IX spi_sdo__i8 (.D(spi_sdo_39__N_145[8]), .SP(clk_enable_961), 
            .CD(n30185), .CK(clk), .Q(spi_sdo[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i8.GSR = "DISABLED";
    FD1P3AX spi_sdo_r__i2 (.D(n23426), .SP(clk_enable_963), .CK(clk), 
            .Q(spi_sdo_r[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i2.GSR = "DISABLED";
    FD1P3IX spi_sdo__i9 (.D(spi_sdo_39__N_145[9]), .SP(clk_enable_961), 
            .CD(n30185), .CK(clk), .Q(spi_sdo[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i9.GSR = "DISABLED";
    FD1P3AX spi_sdo_r__i3 (.D(n23430), .SP(clk_enable_963), .CK(clk), 
            .Q(spi_sdo_r[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i3.GSR = "DISABLED";
    FD1P3IX spi_sdo__i2 (.D(spi_sdo_39__N_145[2]), .SP(clk_enable_961), 
            .CD(n30185), .CK(clk), .Q(spi_sdo[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i2.GSR = "DISABLED";
    FD1P3AX spi_sdo_r__i1 (.D(n23423), .SP(clk_enable_963), .CK(clk), 
            .Q(spi_sdo_r[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i1.GSR = "DISABLED";
    FD1P3AX spi_sdo_r__i4 (.D(n23428), .SP(clk_enable_963), .CK(clk), 
            .Q(spi_sdo_r[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=177, LSE_RLINE=197 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i4.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_806 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[0]), 
         .Z(n23424)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_806.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_807 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[7]), 
         .Z(n23427)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_807.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_808 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[5]), 
         .Z(n23429)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_808.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_809 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[6]), 
         .Z(n23425)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_809.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_810 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[2]), 
         .Z(n23426)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_810.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_811 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[3]), 
         .Z(n23430)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_811.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_812 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[1]), 
         .Z(n23423)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_812.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_813 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[4]), 
         .Z(n23428)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_813.init = 16'h8080;
    LUT4 i23636_2_lut_rep_739 (.A(spi_addr_r[1]), .B(spi_addr_r[4]), .Z(n30139)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23636_2_lut_rep_739.init = 16'heeee;
    LUT4 i23746_2_lut_3_lut (.A(spi_addr_r[1]), .B(spi_addr_r[4]), .C(spi_addr_r[0]), 
         .Z(n28448)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i23746_2_lut_3_lut.init = 16'hfefe;
    LUT4 i23690_2_lut_rep_740 (.A(spi_addr_r[6]), .B(spi_addr_r[7]), .Z(n30140)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23690_2_lut_rep_740.init = 16'heeee;
    LUT4 i23790_3_lut_4_lut (.A(spi_addr_r[6]), .B(spi_addr_r[7]), .C(spi_addr_r[5]), 
         .D(spi_cmd_r[2]), .Z(n28492)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23790_3_lut_4_lut.init = 16'hfffe;
    LUT4 i23786_2_lut_3_lut (.A(spi_addr_r[6]), .B(spi_addr_r[7]), .C(spi_addr_r[0]), 
         .Z(n28488)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i23786_2_lut_3_lut.init = 16'hfefe;
    LUT4 i23680_2_lut_rep_741 (.A(spi_addr_r[3]), .B(spi_addr_r[1]), .Z(n30141)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23680_2_lut_rep_741.init = 16'heeee;
    LUT4 i23796_2_lut_3_lut_4_lut (.A(spi_addr_r[3]), .B(spi_addr_r[1]), 
         .C(spi_addr_r[2]), .D(n30144), .Z(n28498)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23796_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i23824_3_lut_4_lut (.A(spi_addr_r[3]), .B(spi_addr_r[1]), .C(spi_addr_r[2]), 
         .D(n28384), .Z(n28526)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23824_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_742 (.A(spi_cmd_r[4]), .B(spi_cmd_r[5]), .Z(n30142)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_742.init = 16'h8888;
    LUT4 i1_2_lut_rep_644_3_lut (.A(spi_cmd_r[4]), .B(spi_cmd_r[5]), .C(spi_cmd_r[1]), 
         .Z(n30044)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_644_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_814 (.A(spi_cmd_r[4]), .B(spi_cmd_r[5]), .C(spi_addr_r[0]), 
         .Z(n25643)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_3_lut_adj_814.init = 16'h8080;
    LUT4 i1_2_lut_rep_611_3_lut_4_lut (.A(spi_cmd_r[4]), .B(spi_cmd_r[5]), 
         .C(spi_cmd_r[3]), .D(spi_cmd_r[1]), .Z(n30011)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_611_3_lut_4_lut.init = 16'h0800;
    LUT4 i1_2_lut_rep_616_3_lut_4_lut (.A(spi_cmd_r[4]), .B(spi_cmd_r[5]), 
         .C(spi_cmd_r[3]), .D(spi_cmd_r[1]), .Z(n30016)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_616_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_664_3_lut (.A(spi_cmd_r[4]), .B(spi_cmd_r[5]), .C(spi_cmd_r[1]), 
         .Z(n30064)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_664_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_rep_636_3_lut_4_lut (.A(spi_cmd_r[4]), .B(spi_cmd_r[5]), 
         .C(spi_cmd_r[3]), .D(spi_cmd_r[1]), .Z(n30036)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_636_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_815 (.A(spi_cmd_r[4]), .B(spi_cmd_r[5]), 
         .C(spi_cmd_r[3]), .D(spi_cmd_r[1]), .Z(n23537)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_3_lut_4_lut_adj_815.init = 16'h0008;
    LUT4 i23610_2_lut_rep_744 (.A(spi_addr_r[4]), .B(spi_addr_r[6]), .Z(n30144)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23610_2_lut_rep_744.init = 16'heeee;
    LUT4 i23800_3_lut_rep_670_4_lut (.A(spi_addr_r[4]), .B(spi_addr_r[6]), 
         .C(spi_addr_r[2]), .D(n30155), .Z(n30070)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23800_3_lut_rep_670_4_lut.init = 16'hfffe;
    LUT4 i23582_2_lut_rep_750 (.A(spi_addr_r[2]), .B(spi_addr_r[3]), .Z(n30150)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23582_2_lut_rep_750.init = 16'heeee;
    LUT4 i23792_2_lut_3_lut_4_lut (.A(spi_addr_r[2]), .B(spi_addr_r[3]), 
         .C(n30213), .D(n30214), .Z(n28494)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23792_2_lut_3_lut_4_lut.init = 16'hfffe;
    wb_ctrl wb_ctrl_inst (.wb_cyc_i(wb_cyc_i), .clk(clk), .clk_enable_172(clk_enable_172), 
            .\wb_adr_i[0] (wb_adr_i[0]), .\address[0] (address[0]), .wb_we_i(wb_we_i), 
            .wb_we_i_N_344(wb_we_i_N_344), .wb_dat_i({wb_dat_i}), .wr_data({wr_data}), 
            .wb_sm(wb_sm), .spi_cmd_start(spi_cmd_start), .\address_7__N_549[1] (address_7__N_549[1]), 
            .\address_7__N_565[1] (address_7__N_565[1]), .wr_en(wr_en), 
            .wr_en_N_355(wr_en_N_355), .\wb_adr_i[1] (wb_adr_i[1]), .\address[1] (address[1]), 
            .\wb_adr_i[6] (wb_adr_i[6]), .n31069(n31069), .rd_en(rd_en), 
            .n29(n29)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/spi_slave_top.v(179[12] 196[15])
    spi_slave_efb spi_slave_efb_inst (.clk(clk), .n30185(n30185), .wb_cyc_i(wb_cyc_i), 
            .wb_we_i(wb_we_i), .GND_net(GND_net), .\wb_adr_i[6] (wb_adr_i[6]), 
            .\wb_adr_i[1] (wb_adr_i[1]), .\wb_adr_i[0] (wb_adr_i[0]), .wb_dat_i({wb_dat_i}), 
            .spi_scsn_c(spi_scsn_c), .wb_dat_o({wb_dat_o}), .\address_7__N_549[1] (address_7__N_549[1]), 
            .spi_mosi_oe(spi_mosi_oe), .spi_mosi_o(spi_mosi_o), .spi_miso_oe(spi_miso_oe), 
            .spi_miso_o(spi_miso_o), .spi_clk_oe(spi_clk_oe), .spi_clk_o(spi_clk_o), 
            .spi_mosi_i(spi_mosi_i), .spi_miso_i(spi_miso_i), .spi_clk_i(spi_clk_i), 
            .VCC_net(VCC_net), .wb_sm(wb_sm), .clk_enable_172(clk_enable_172)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/s_links/sources/spi_slave_top.v(162[18] 176[15])
    spi_ctrl spi_ctrl_inst (.quad_buffer({quad_buffer}), .quad_count({quad_count}), 
            .\spi_data_out_r_39__N_1083[31] (\spi_data_out_r_39__N_1083[31] ), 
            .spi_addr({spi_addr}), .spi_cmd({spi_cmd[15:3], \spi_cmd[2] , 
            spi_cmd[1:0]}), .clk(clk), .\spi_data[0] (spi_data[0]), .wb_dat_o({wb_dat_o}), 
            .\spi_data_out_r_39__N_1083[29] (\spi_data_out_r_39__N_1083[29] ), 
            .wr_en_N_355(wr_en_N_355), .wr_data({wr_data}), .\address[0] (address[0]), 
            .rd_en(rd_en), .wr_en(wr_en), .spi_scsn_c(spi_scsn_c), .\address_7__N_549[1] (address_7__N_549[1]), 
            .\spi_data_out_r_39__N_1083[19] (\spi_data_out_r_39__N_1083[19] ), 
            .\spi_data_out_r_39__N_1083[18] (\spi_data_out_r_39__N_1083[18] ), 
            .quad_buffer_adj_321({quad_buffer_adj_644}), .quad_count_adj_322({quad_count_adj_645}), 
            .\spi_data_out_r_39__N_2023[26] (\spi_data_out_r_39__N_2023[26] ), 
            .n30198(n30198), .n32(n32), .clear_intrpt_N_2717(clear_intrpt_N_2717), 
            .\address_7__N_565[1] (address_7__N_565[1]), .resetn_c(resetn_c), 
            .spi_addr_valid(spi_addr_valid), .n47(n47), .clear_intrpt_N_2930(clear_intrpt_N_2930), 
            .clear_intrpt_N_2788(clear_intrpt_N_2788), .clear_intrpt_N_2859(clear_intrpt_N_2859), 
            .n47_adj_74(n47_adj_400), .quad_buffer_adj_323({quad_buffer_adj_646}), 
            .quad_count_adj_324({quad_count_adj_647}), .\spi_data_out_r_39__N_2493[29] (\spi_data_out_r_39__N_2493[29] ), 
            .\spi_data_out_r_39__N_2493[28] (\spi_data_out_r_39__N_2493[28] ), 
            .\spi_data_out_r_39__N_2493[27] (\spi_data_out_r_39__N_2493[27] ), 
            .\spi_data_out_r_39__N_2493[26] (\spi_data_out_r_39__N_2493[26] ), 
            .n29997(n29997), .n29991(n29991), .\spi_data_out_r_39__N_2493[25] (\spi_data_out_r_39__N_2493[25] ), 
            .\spi_data_out_r_39__N_2493[24] (\spi_data_out_r_39__N_2493[24] ), 
            .\spi_data_out_r_39__N_2493[23] (\spi_data_out_r_39__N_2493[23] ), 
            .\spi_data_out_r_39__N_2493[22] (\spi_data_out_r_39__N_2493[22] ), 
            .\spi_data_out_r_39__N_2493[21] (\spi_data_out_r_39__N_2493[21] ), 
            .\spi_data_out_r_39__N_2493[20] (\spi_data_out_r_39__N_2493[20] ), 
            .\spi_data_out_r_39__N_2493[19] (\spi_data_out_r_39__N_2493[19] ), 
            .\spi_data[31] (spi_data[31]), .\spi_data_out_r_39__N_2493[18] (\spi_data_out_r_39__N_2493[18] ), 
            .\spi_data_out_r_39__N_2493[17] (\spi_data_out_r_39__N_2493[17] ), 
            .\spi_data_out_r_39__N_2493[16] (\spi_data_out_r_39__N_2493[16] ), 
            .\spi_data_out_r_39__N_2493[15] (\spi_data_out_r_39__N_2493[15] ), 
            .\spi_data_out_r_39__N_2493[14] (\spi_data_out_r_39__N_2493[14] ), 
            .\spi_data_out_r_39__N_2493[13] (\spi_data_out_r_39__N_2493[13] ), 
            .\spi_data_out_r_39__N_2493[12] (\spi_data_out_r_39__N_2493[12] ), 
            .\spi_data_out_r_39__N_2493[11] (\spi_data_out_r_39__N_2493[11] ), 
            .\spi_data_out_r_39__N_2493[10] (\spi_data_out_r_39__N_2493[10] ), 
            .\spi_data[30] (spi_data[30]), .\spi_data[29] (spi_data[29]), 
            .\spi_data[28] (spi_data[28]), .\spi_data[27] (spi_data[27]), 
            .\spi_data[26] (spi_data[26]), .\spi_data[25] (spi_data[25]), 
            .\spi_data[24] (spi_data[24]), .\spi_data[23] (spi_data[23]), 
            .\spi_data[22] (spi_data[22]), .\spi_data_out_r_39__N_2493[9] (\spi_data_out_r_39__N_2493[9] ), 
            .\spi_data_out_r_39__N_2493[8] (\spi_data_out_r_39__N_2493[8] ), 
            .\spi_data[21] (spi_data[21]), .\spi_data[20] (spi_data[20]), 
            .\spi_data[19] (spi_data[19]), .\spi_data[18] (spi_data[18]), 
            .\spi_data[17] (spi_data[17]), .\spi_data_out_r_39__N_2493[7] (\spi_data_out_r_39__N_2493[7] ), 
            .\spi_data[16] (spi_data[16]), .\spi_data[15] (spi_data[15]), 
            .\spi_data[14] (spi_data[14]), .\spi_data[13] (spi_data[13]), 
            .\spi_data[12] (spi_data[12]), .\spi_data[11] (spi_data[11]), 
            .\spi_data[10] (spi_data[10]), .\spi_data[9] (spi_data[9]), 
            .\spi_data[8] (spi_data[8]), .\spi_data[7] (spi_data[7]), .\spi_data[6] (spi_data[6]), 
            .\spi_data[5] (spi_data[5]), .\spi_data[4] (spi_data[4]), .\spi_data[3] (spi_data[3]), 
            .\spi_data_out_r_39__N_1083[9] (\spi_data_out_r_39__N_1083[9] ), 
            .\spi_data[2] (spi_data[2]), .\spi_data[1] (spi_data[1]), .\spi_data_out_r_39__N_1083[8] (\spi_data_out_r_39__N_1083[8] ), 
            .\spi_data_out_r_39__N_2493[6] (\spi_data_out_r_39__N_2493[6] ), 
            .\spi_data_out_r_39__N_2493[5] (\spi_data_out_r_39__N_2493[5] ), 
            .\spi_data_out_r_39__N_2493[4] (\spi_data_out_r_39__N_2493[4] ), 
            .\spi_data_out_r_39__N_2493[3] (\spi_data_out_r_39__N_2493[3] ), 
            .\spi_data_out_r_39__N_2493[2] (\spi_data_out_r_39__N_2493[2] ), 
            .\spi_data_out_r_39__N_2493[1] (\spi_data_out_r_39__N_2493[1] ), 
            .\spi_data_out_r_39__N_2023[20] (\spi_data_out_r_39__N_2023[20] ), 
            .quad_buffer_adj_325({quad_buffer_adj_648}), .quad_count_adj_326({quad_count_adj_649}), 
            .\spi_data_out_r_39__N_2258[0] (\spi_data_out_r_39__N_2258[0] ), 
            .\spi_data_out_r_39__N_2258[31] (\spi_data_out_r_39__N_2258[31] ), 
            .\spi_data_out_r_39__N_2258[30] (\spi_data_out_r_39__N_2258[30] ), 
            .\spi_data_out_r_39__N_2258[29] (\spi_data_out_r_39__N_2258[29] ), 
            .\spi_data_out_r_39__N_2258[28] (\spi_data_out_r_39__N_2258[28] ), 
            .\spi_data_out_r_39__N_2258[27] (\spi_data_out_r_39__N_2258[27] ), 
            .\spi_data_out_r_39__N_2258[26] (\spi_data_out_r_39__N_2258[26] ), 
            .n26779(n26779), .\spi_data_out_r_39__N_2258[25] (\spi_data_out_r_39__N_2258[25] ), 
            .\spi_data_out_r_39__N_2258[24] (\spi_data_out_r_39__N_2258[24] ), 
            .\spi_data_out_r_39__N_1083[22] (\spi_data_out_r_39__N_1083[22] ), 
            .\spi_data_out_r_39__N_2258[23] (\spi_data_out_r_39__N_2258[23] ), 
            .\spi_data_out_r_39__N_2258[22] (\spi_data_out_r_39__N_2258[22] ), 
            .\spi_data_out_r_39__N_2258[21] (\spi_data_out_r_39__N_2258[21] ), 
            .\spi_data_out_r_39__N_2258[20] (\spi_data_out_r_39__N_2258[20] ), 
            .\spi_data_out_r_39__N_2258[19] (\spi_data_out_r_39__N_2258[19] ), 
            .\spi_data_out_r_39__N_2258[18] (\spi_data_out_r_39__N_2258[18] ), 
            .n47_adj_203(n47_adj_529), .\spi_data_out_r_39__N_2258[17] (\spi_data_out_r_39__N_2258[17] ), 
            .\spi_data_out_r_39__N_2258[16] (\spi_data_out_r_39__N_2258[16] ), 
            .\spi_data_out_r_39__N_2258[15] (\spi_data_out_r_39__N_2258[15] ), 
            .\spi_data_out_r_39__N_2258[14] (\spi_data_out_r_39__N_2258[14] ), 
            .\spi_data_out_r_39__N_2258[13] (\spi_data_out_r_39__N_2258[13] ), 
            .\spi_data_out_r_39__N_2258[12] (\spi_data_out_r_39__N_2258[12] ), 
            .\spi_data_out_r_39__N_2258[11] (\spi_data_out_r_39__N_2258[11] ), 
            .\spi_data_out_r_39__N_2258[10] (\spi_data_out_r_39__N_2258[10] ), 
            .\spi_data_out_r_39__N_2258[9] (\spi_data_out_r_39__N_2258[9] ), 
            .n30019(n30019), .n47_adj_204(n47_adj_530), .\spi_data_out_r_39__N_2258[8] (\spi_data_out_r_39__N_2258[8] ), 
            .\address[1] (address[1]), .\spi_data_out_r_39__N_2258[7] (\spi_data_out_r_39__N_2258[7] ), 
            .n30027(n30027), .n47_adj_205(n47_adj_531), .\spi_data_out_r_39__N_2258[6] (\spi_data_out_r_39__N_2258[6] ), 
            .\spi_data_out_r_39__N_2258[5] (\spi_data_out_r_39__N_2258[5] ), 
            .\spi_data_out_r_39__N_2258[4] (\spi_data_out_r_39__N_2258[4] ), 
            .\spi_data_out_r_39__N_2258[3] (\spi_data_out_r_39__N_2258[3] ), 
            .\spi_data_out_r_39__N_1083[17] (\spi_data_out_r_39__N_1083[17] ), 
            .\spi_data_out_r_39__N_2258[2] (\spi_data_out_r_39__N_2258[2] ), 
            .\spi_data_out_r_39__N_2023[19] (\spi_data_out_r_39__N_2023[19] ), 
            .\spi_data_out_r_39__N_2258[1] (\spi_data_out_r_39__N_2258[1] ), 
            .\SLO_buf[4] (\SLO_buf[4] ), .\SLO_buf[14] (\SLO_buf[14] ), 
            .\spi_data_out_r_39__N_5105[0] (\spi_data_out_r_39__N_5105[0] ), 
            .\SLO_buf[3] (\SLO_buf[3] ), .\SLO_buf[9] (\SLO_buf[9] ), .\spi_data_out_r_39__N_5105[35] (\spi_data_out_r_39__N_5105[35] ), 
            .\SLO_buf[2] (\SLO_buf[2] ), .\SLO_buf[8] (\SLO_buf[8] ), .\spi_data_out_r_39__N_5105[34] (\spi_data_out_r_39__N_5105[34] ), 
            .\SLO_buf[1] (\SLO_buf[1] ), .\SLO_buf[7] (\SLO_buf[7] ), .\spi_data_out_r_39__N_5105[33] (\spi_data_out_r_39__N_5105[33] ), 
            .quad_buffer_adj_327({quad_buffer_adj_650}), .quad_count_adj_328({quad_count_adj_651}), 
            .\spi_data_out_r_39__N_1553[0] (\spi_data_out_r_39__N_1553[0] ), 
            .\spi_data_out_r_39__N_1553[31] (\spi_data_out_r_39__N_1553[31] ), 
            .\SLO_buf[0] (\SLO_buf[0] ), .\SLO_buf[6] (\SLO_buf[6] ), .\spi_data_out_r_39__N_5105[32] (\spi_data_out_r_39__N_5105[32] ), 
            .\SLO_buf[19] (\SLO_buf[19] ), .\SLO_buf[29] (\SLO_buf[29] ), 
            .\spi_data_out_r_39__N_5105[15] (\spi_data_out_r_39__N_5105[15] ), 
            .\spi_data_out_r_39__N_1553[30] (\spi_data_out_r_39__N_1553[30] ), 
            .\spi_data_out_r_39__N_1553[29] (\spi_data_out_r_39__N_1553[29] ), 
            .\spi_data_out_r_39__N_1553[28] (\spi_data_out_r_39__N_1553[28] ), 
            .\spi_data_out_r_39__N_1553[27] (\spi_data_out_r_39__N_1553[27] ), 
            .\SLO_buf[18] (\SLO_buf[18] ), .\SLO_buf[28] (\SLO_buf[28] ), 
            .\spi_data_out_r_39__N_5105[14] (\spi_data_out_r_39__N_5105[14] ), 
            .\spi_data_out_r_39__N_1553[26] (\spi_data_out_r_39__N_1553[26] ), 
            .\SLO_buf[17] (\SLO_buf[17] ), .\SLO_buf[27] (\SLO_buf[27] ), 
            .\spi_data_out_r_39__N_5105[13] (\spi_data_out_r_39__N_5105[13] ), 
            .\spi_data_out_r_39__N_2023[25] (\spi_data_out_r_39__N_2023[25] ), 
            .\spi_data_out_r_39__N_1553[25] (\spi_data_out_r_39__N_1553[25] ), 
            .\spi_data_out_r_39__N_1553[24] (\spi_data_out_r_39__N_1553[24] ), 
            .wb_sm(wb_sm), .wb_we_i_N_344(wb_we_i_N_344), .\SLO_buf[16] (\SLO_buf[16] ), 
            .\SLO_buf[26] (\SLO_buf[26] ), .\spi_data_out_r_39__N_5105[12] (\spi_data_out_r_39__N_5105[12] ), 
            .\spi_data_out_r_39__N_1553[23] (\spi_data_out_r_39__N_1553[23] ), 
            .\SLO_buf[15] (\SLO_buf[15] ), .\SLO_buf[25] (\SLO_buf[25] ), 
            .\spi_data_out_r_39__N_5105[11] (\spi_data_out_r_39__N_5105[11] ), 
            .\SLO_buf[24] (\SLO_buf[24] ), .\spi_data_out_r_39__N_5105[10] (\spi_data_out_r_39__N_5105[10] ), 
            .\spi_data_out_r_39__N_1553[22] (\spi_data_out_r_39__N_1553[22] ), 
            .\SLO_buf[13] (\SLO_buf[13] ), .\SLO_buf[23] (\SLO_buf[23] ), 
            .\spi_data_out_r_39__N_5105[9] (\spi_data_out_r_39__N_5105[9] ), 
            .\spi_data_out_r_39__N_1553[21] (\spi_data_out_r_39__N_1553[21] ), 
            .\spi_data_out_r_39__N_1553[20] (\spi_data_out_r_39__N_1553[20] ), 
            .\spi_data_out_r_39__N_1553[19] (\spi_data_out_r_39__N_1553[19] ), 
            .\spi_data_out_r_39__N_1553[18] (\spi_data_out_r_39__N_1553[18] ), 
            .\spi_data_out_r_39__N_1553[17] (\spi_data_out_r_39__N_1553[17] ), 
            .\spi_data_out_r_39__N_1553[16] (\spi_data_out_r_39__N_1553[16] ), 
            .\spi_data_out_r_39__N_1083[16] (\spi_data_out_r_39__N_1083[16] ), 
            .\spi_data_out_r_39__N_1553[15] (\spi_data_out_r_39__N_1553[15] ), 
            .\spi_data_out_r_39__N_1553[14] (\spi_data_out_r_39__N_1553[14] ), 
            .\spi_data_out_r_39__N_1553[13] (\spi_data_out_r_39__N_1553[13] ), 
            .\spi_data_out_r_39__N_1083[15] (\spi_data_out_r_39__N_1083[15] ), 
            .GND_net(GND_net), .\SLO_buf[12] (\SLO_buf[12] ), .\SLO_buf[22] (\SLO_buf[22] ), 
            .\spi_data_out_r_39__N_5105[8] (\spi_data_out_r_39__N_5105[8] ), 
            .\spi_data_out_r_39__N_1553[12] (\spi_data_out_r_39__N_1553[12] ), 
            .\SLO_buf[11] (\SLO_buf[11] ), .\SLO_buf[21] (\SLO_buf[21] ), 
            .\spi_data_out_r_39__N_5105[7] (\spi_data_out_r_39__N_5105[7] ), 
            .\spi_data_out_r_39__N_1553[11] (\spi_data_out_r_39__N_1553[11] ), 
            .\SLO_buf[10] (\SLO_buf[10] ), .\SLO_buf[20] (\SLO_buf[20] ), 
            .\spi_data_out_r_39__N_5105[6] (\spi_data_out_r_39__N_5105[6] ), 
            .\spi_data_out_r_39__N_5105[5] (\spi_data_out_r_39__N_5105[5] ), 
            .\spi_data_out_r_39__N_1553[10] (\spi_data_out_r_39__N_1553[10] ), 
            .\spi_data_out_r_39__N_5105[4] (\spi_data_out_r_39__N_5105[4] ), 
            .\spi_data_out_r_39__N_1553[9] (\spi_data_out_r_39__N_1553[9] ), 
            .\spi_data_out_r_39__N_1553[8] (\spi_data_out_r_39__N_1553[8] ), 
            .\spi_data_out_r_39__N_1553[7] (\spi_data_out_r_39__N_1553[7] ), 
            .\spi_data_out_r_39__N_1553[6] (\spi_data_out_r_39__N_1553[6] ), 
            .\spi_data_out_r_39__N_5105[3] (\spi_data_out_r_39__N_5105[3] ), 
            .\spi_data_out_r_39__N_1553[5] (\spi_data_out_r_39__N_1553[5] ), 
            .\spi_data_out_r_39__N_1553[4] (\spi_data_out_r_39__N_1553[4] ), 
            .\spi_data_out_r_39__N_1553[3] (\spi_data_out_r_39__N_1553[3] ), 
            .\spi_data_out_r_39__N_2023[18] (\spi_data_out_r_39__N_2023[18] ), 
            .\spi_data_out_r_39__N_1553[2] (\spi_data_out_r_39__N_1553[2] ), 
            .\spi_data_out_r_39__N_1553[1] (\spi_data_out_r_39__N_1553[1] ), 
            .n47_adj_270(n47_adj_596), .spi_cmd_start(spi_cmd_start), .\spi_data_out_r_39__N_5105[2] (\spi_data_out_r_39__N_5105[2] ), 
            .\SLO_buf[5] (\SLO_buf[5] ), .\spi_data_out_r_39__N_5105[1] (\spi_data_out_r_39__N_5105[1] ), 
            .n29(n29), .spi_data_out_r_39__N_2338(spi_data_out_r_39__N_2338), 
            .n47_adj_271(n47_adj_597), .\spi_data_out_r_39__N_1083[14] (\spi_data_out_r_39__N_1083[14] ), 
            .\spi_data_out_r_39__N_1083[13] (\spi_data_out_r_39__N_1083[13] ), 
            .n30102(n30102), .\SLO_buf[4]_adj_272 (\SLO_buf[4]_adj_598 ), 
            .\SLO_buf[14]_adj_273 (\SLO_buf[14]_adj_599 ), .\spi_data_out_r_39__N_4419[0] (\spi_data_out_r_39__N_4419[0] ), 
            .mem_rdata({mem_rdata}), .\SLO_buf[3]_adj_274 (\SLO_buf[3]_adj_600 ), 
            .\SLO_buf[9]_adj_275 (\SLO_buf[9]_adj_601 ), .\spi_data_out_r_39__N_4419[35] (\spi_data_out_r_39__N_4419[35] ), 
            .spi_data_out_r_39__N_4505(spi_data_out_r_39__N_4505), .\spi_data_out_r_39__N_2023[17] (\spi_data_out_r_39__N_2023[17] ), 
            .\spi_data_out_r_39__N_2023[16] (\spi_data_out_r_39__N_2023[16] ), 
            .\spi_data_out_r_39__N_1083[7] (\spi_data_out_r_39__N_1083[7] ), 
            .\spi_data_out_r_39__N_1083[6] (\spi_data_out_r_39__N_1083[6] ), 
            .\spi_data_out_r_39__N_1083[20] (\spi_data_out_r_39__N_1083[20] ), 
            .\spi_data_out_r_39__N_2023[15] (\spi_data_out_r_39__N_2023[15] ), 
            .\status_cntr[12] (\status_cntr[12] ), .n25212(n25212), .\SLO_buf[2]_adj_276 (\SLO_buf[2]_adj_602 ), 
            .\SLO_buf[8]_adj_277 (\SLO_buf[8]_adj_603 ), .\spi_data_out_r_39__N_4419[34] (\spi_data_out_r_39__N_4419[34] ), 
            .\spi_data_out_r_39__N_2023[14] (\spi_data_out_r_39__N_2023[14] ), 
            .\SLO_buf[1]_adj_278 (\SLO_buf[1]_adj_604 ), .\SLO_buf[7]_adj_279 (\SLO_buf[7]_adj_605 ), 
            .\spi_data_out_r_39__N_4419[33] (\spi_data_out_r_39__N_4419[33] ), 
            .\SLO_buf[0]_adj_280 (\SLO_buf[0]_adj_606 ), .\SLO_buf[6]_adj_281 (\SLO_buf[6]_adj_607 ), 
            .\spi_data_out_r_39__N_4419[32] (\spi_data_out_r_39__N_4419[32] ), 
            .clear_intrpt_N_3072(clear_intrpt_N_3072), .\spi_data_out_r_39__N_2023[13] (\spi_data_out_r_39__N_2023[13] ), 
            .\SLO_buf[19]_adj_282 (\SLO_buf[19]_adj_608 ), .\SLO_buf[29]_adj_283 (\SLO_buf[29]_adj_609 ), 
            .\spi_data_out_r_39__N_4419[15] (\spi_data_out_r_39__N_4419[15] ), 
            .\spi_data_out_r_39__N_1083[5] (\spi_data_out_r_39__N_1083[5] ), 
            .\spi_data_out_r_39__N_1083[4] (\spi_data_out_r_39__N_1083[4] ), 
            .\spi_data_out_r_39__N_2023[12] (\spi_data_out_r_39__N_2023[12] ), 
            .\SLO_buf[18]_adj_284 (\SLO_buf[18]_adj_610 ), .\SLO_buf[28]_adj_285 (\SLO_buf[28]_adj_611 ), 
            .\spi_data_out_r_39__N_4419[14] (\spi_data_out_r_39__N_4419[14] ), 
            .\SLO_buf[17]_adj_286 (\SLO_buf[17]_adj_612 ), .\SLO_buf[27]_adj_287 (\SLO_buf[27]_adj_613 ), 
            .\spi_data_out_r_39__N_4419[13] (\spi_data_out_r_39__N_4419[13] ), 
            .\spi_data_out_r_39__N_1083[12] (\spi_data_out_r_39__N_1083[12] ), 
            .spi_data_out_r_39__N_4848(spi_data_out_r_39__N_4848), .\spi_data_out_r_39__N_1083[3] (\spi_data_out_r_39__N_1083[3] ), 
            .\spi_data_out_r_39__N_1083[2] (\spi_data_out_r_39__N_1083[2] ), 
            .\spi_data_out_r_39__N_2023[11] (\spi_data_out_r_39__N_2023[11] ), 
            .\SLO_buf[16]_adj_288 (\SLO_buf[16]_adj_614 ), .\SLO_buf[26]_adj_289 (\SLO_buf[26]_adj_615 ), 
            .\spi_data_out_r_39__N_4419[12] (\spi_data_out_r_39__N_4419[12] ), 
            .\spi_data_out_r_39__N_2023[10] (\spi_data_out_r_39__N_2023[10] ), 
            .\SLO_buf[15]_adj_290 (\SLO_buf[15]_adj_616 ), .\SLO_buf[25]_adj_291 (\SLO_buf[25]_adj_617 ), 
            .\spi_data_out_r_39__N_4419[11] (\spi_data_out_r_39__N_4419[11] ), 
            .\SLO_buf[24]_adj_292 (\SLO_buf[24]_adj_618 ), .\spi_data_out_r_39__N_4419[10] (\spi_data_out_r_39__N_4419[10] ), 
            .\SLO_buf[13]_adj_293 (\SLO_buf[13]_adj_619 ), .\SLO_buf[23]_adj_294 (\SLO_buf[23]_adj_620 ), 
            .\spi_data_out_r_39__N_4419[9] (\spi_data_out_r_39__N_4419[9] ), 
            .\SLO_buf[12]_adj_295 (\SLO_buf[12]_adj_621 ), .\SLO_buf[22]_adj_296 (\SLO_buf[22]_adj_622 ), 
            .\spi_data_out_r_39__N_4419[8] (\spi_data_out_r_39__N_4419[8] ), 
            .n30185(n30185), .n25885(n25885), .n30087(n30087), .\quad_homing[1] (\quad_homing[1] ), 
            .n1(n1), .spi_sdo_valid(spi_sdo_valid), .clk_enable_963(clk_enable_963), 
            .n30010(n30010), .\spi_addr_r[0] (spi_addr_r[0]), .clk_enable_686(clk_enable_686), 
            .spi_cmd_valid(spi_cmd_valid), .spi_scsn_dly(spi_scsn_dly), 
            .clk_enable_776(clk_enable_776), .n26077(n26077), .n24066(n24066), 
            .n30062(n30062), .clk_enable_260(clk_enable_260), .clear_intrpt(clear_intrpt_adj_623), 
            .intrpt_out_N_2642(intrpt_out_N_2642), .clear_intrpt_adj_297(clear_intrpt_adj_333), 
            .intrpt_out_N_3068(intrpt_out_N_3068), .n28540(n28540), .n30035(n30035), 
            .n23537(n23537), .clk_enable_263(clk_enable_263), .quad_set_valid_N_1158(quad_set_valid_N_1158), 
            .clk_enable_807(clk_enable_807), .n20598(n20598), .n8400(n8400), 
            .n12467(n12467), .n20647(n20647), .n18654(n18654), .n12435(n12435), 
            .n4(n4), .n30070(n30070), .n26873(n26873), .clk_enable_320(clk_enable_320), 
            .n25877(n25877), .n30075(n30075), .\quad_homing[1]_adj_298 (\quad_homing[1]_adj_624 ), 
            .n1_adj_299(n1_adj_625), .n30199(n30199), .n23916(n23916), 
            .n26821(n26821), .clk_enable_684(clk_enable_684), .n26089(n26089), 
            .n26091(n26091), .clk_enable_255(clk_enable_255), .EM_STOP(EM_STOP), 
            .clk_enable_259(clk_enable_259), .n29996(n29996), .clk_enable_23(clk_enable_23), 
            .n26947(n26947), .clk_enable_253(clk_enable_253), .pwm_out_N_3169(pwm_out_N_3169), 
            .pwm_out_N_3153(pwm_out_N_3153), .clk_enable_15(clk_enable_15), 
            .\spi_addr_r[7] (spi_addr_r[7]), .n26107(n26107), .n30214(n30214), 
            .n26113(n26113), .clear_intrpt_adj_300(clear_intrpt_adj_626), 
            .intrpt_out_N_2997(intrpt_out_N_2997), .n25993(n25993), .clk_enable_687(clk_enable_687), 
            .n30045(n30045), .n28524(n28524), .clk_enable_759(clk_enable_759), 
            .clk_enable_48(clk_enable_48), .clk_enable_624(clk_enable_624), 
            .n30033(n30033), .n23526(n23526), .clk_enable_727(clk_enable_727), 
            .n11008(n11008), .pwm_out_1_N_6491(pwm_out_1_N_6491), .clk_enable_613(clk_enable_613), 
            .spi_sdo_valid_N_296(spi_sdo_valid_N_296), .clk_enable_961(clk_enable_961), 
            .n30011(n30011), .n26957(n26957), .clk_enable_520(clk_enable_520), 
            .n28364(n28364), .n24065(n24065), .n26033(n26033), .clk_enable_232(clk_enable_232), 
            .clk_enable_254(clk_enable_254), .n29995(n29995), .clk_enable_28(clk_enable_28), 
            .n28514(n28514), .n26563(n26563), .clk_enable_226(clk_enable_226), 
            .clk_enable_639(clk_enable_639), .clk_enable_228(clk_enable_228), 
            .pwm_out_3_N_6530(pwm_out_3_N_6530), .clk_enable_1105(clk_enable_1105), 
            .pwm_out_4_N_6549(pwm_out_4_N_6549), .clk_enable_1107(clk_enable_1107), 
            .n26841(n26841), .n26843(n26843), .clk_enable_757(clk_enable_757), 
            .n26023(n26023), .n28366(n28366), .clk_enable_245(clk_enable_245), 
            .pwm_out_2_N_6511(pwm_out_2_N_6511), .clk_enable_22(clk_enable_22), 
            .n30022(n30022), .n26415(n26415), .clk_enable_488(clk_enable_488), 
            .n26633(n26633), .clk_enable_641(clk_enable_641), .n25833(n25833), 
            .clk_enable_638(clk_enable_638), .n30036(n30036), .n26435(n26435), 
            .clk_enable_959(clk_enable_959), .n18440(n18440), .n26249(n26249), 
            .clk_enable_235(clk_enable_235), .clear_intrpt_adj_301(clear_intrpt_adj_335), 
            .intrpt_out_N_2713(intrpt_out_N_2713), .n57(n57), .reset_r_N_4129(reset_r_N_4129), 
            .clk_enable_761(clk_enable_761), .n30080(n30080), .n29998(n29998), 
            .n26539(n26539), .clk_enable_738(clk_enable_738), .n25881(n25881), 
            .n30095(n30095), .\quad_homing[1]_adj_302 (\quad_homing[1]_adj_627 ), 
            .n1_adj_303(n1_adj_628), .n28516(n28516), .n26515(n26515), 
            .clk_enable_652(clk_enable_652), .quad_set_valid_N_2098(quad_set_valid_N_2098), 
            .clk_enable_683(clk_enable_683), .clk_enable_211(clk_enable_211), 
            .n2109(n2109), .n25893(n25893), .n30055(n30055), .\quad_homing[1]_adj_304 (\quad_homing[1]_adj_629 ), 
            .n1_adj_305(n1_adj_630), .n25869(n25869), .n30043(n30043), 
            .\quad_homing[1]_adj_306 (\quad_homing[1]_adj_631 ), .n1_adj_307(n1_adj_632), 
            .n25873(n25873), .n30091(n30091), .\quad_homing[1]_adj_308 (\quad_homing[1]_adj_633 ), 
            .n1_adj_309(n1_adj_634), .n28476(n28476), .n26059(n26059), 
            .clk_enable_32(clk_enable_32), .clear_intrpt_adj_310(clear_intrpt_adj_334), 
            .intrpt_out_N_2855(intrpt_out_N_2855), .clk_enable_178(clk_enable_178), 
            .clear_intrpt_adj_311(clear_intrpt_adj_332), .intrpt_out_N_2784(intrpt_out_N_2784), 
            .quad_set_valid_N_1393(quad_set_valid_N_1393), .clk_enable_842(clk_enable_842), 
            .n27013(n27013), .clk_enable_627(clk_enable_627), .n26233(n26233), 
            .clk_enable_234(clk_enable_234), .quad_set_valid_N_2333(quad_set_valid_N_2333), 
            .clk_enable_315(clk_enable_315), .\SLO_buf[11]_adj_312 (\SLO_buf[11]_adj_635 ), 
            .\SLO_buf[21]_adj_313 (\SLO_buf[21]_adj_636 ), .\spi_data_out_r_39__N_4419[7] (\spi_data_out_r_39__N_4419[7] ), 
            .clk_enable_256(clk_enable_256), .n29999(n29999), .clk_enable_12(clk_enable_12), 
            .n26587(n26587), .clk_enable_749(clk_enable_749), .clk_enable_388(clk_enable_388), 
            .n26207(n26207), .clk_enable_898(clk_enable_898), .clk_enable_180(clk_enable_180), 
            .n18(n18_adj_637), .n2193(n2193), .\SLO_buf[10]_adj_314 (\SLO_buf[10]_adj_638 ), 
            .\SLO_buf[20]_adj_315 (\SLO_buf[20]_adj_639 ), .\spi_data_out_r_39__N_4419[6] (\spi_data_out_r_39__N_4419[6] ), 
            .clk_enable_244(clk_enable_244), .clear_intrpt_adj_316(clear_intrpt), 
            .intrpt_out_N_2926(intrpt_out_N_2926), .pwm_out_1_N_6306(pwm_out_1_N_6306), 
            .clk_100k_enable_1(clk_100k_enable_1), .n25889(n25889), .n30083(n30083), 
            .\quad_homing[1]_adj_317 (\quad_homing[1]_adj_640 ), .n1_adj_318(n1_adj_641), 
            .clk_enable_595(clk_enable_595), .n30039(n30039), .\spi_data_out_r_39__N_2023[9] (\spi_data_out_r_39__N_2023[9] ), 
            .\spi_data_out_r_39__N_1083[24] (\spi_data_out_r_39__N_1083[24] ), 
            .clear_intrpt_N_3001(clear_intrpt_N_3001), .\spi_data_out_r_39__N_2023[8] (\spi_data_out_r_39__N_2023[8] ), 
            .\spi_data_out_r_39__N_1083[11] (\spi_data_out_r_39__N_1083[11] ), 
            .\spi_data_out_r_39__N_2023[7] (\spi_data_out_r_39__N_2023[7] ), 
            .\spi_data_out_r_39__N_1083[27] (\spi_data_out_r_39__N_1083[27] ), 
            .\spi_data_out_r_39__N_4419[5] (\spi_data_out_r_39__N_4419[5] ), 
            .\spi_data_out_r_39__N_4419[4] (\spi_data_out_r_39__N_4419[4] ), 
            .\spi_data_out_r_39__N_2023[6] (\spi_data_out_r_39__N_2023[6] ), 
            .n27095(n27095), .spi_data_out_r_39__N_1868(spi_data_out_r_39__N_1868), 
            .n29992(n29992), .\spi_data_out_r_39__N_4419[3] (\spi_data_out_r_39__N_4419[3] ), 
            .\spi_data_out_r_39__N_2023[5] (\spi_data_out_r_39__N_2023[5] ), 
            .\spi_data_out_r_39__N_2023[24] (\spi_data_out_r_39__N_2023[24] ), 
            .\spi_data_out_r_39__N_4419[2] (\spi_data_out_r_39__N_4419[2] ), 
            .n28452(n28452), .spi_data_out_r_39__N_5191(spi_data_out_r_39__N_5191), 
            .spi_data_out_r_39__N_5534(spi_data_out_r_39__N_5534), .spi_data_out_r_39__N_5877(spi_data_out_r_39__N_5877), 
            .\spi_data_out_r_39__N_1083[23] (\spi_data_out_r_39__N_1083[23] ), 
            .spi_data_out_r_39__N_6220(spi_data_out_r_39__N_6220), .\spi_data_out_r_39__N_2023[4] (\spi_data_out_r_39__N_2023[4] ), 
            .\spi_data_out_r_39__N_2023[23] (\spi_data_out_r_39__N_2023[23] ), 
            .\spi_data_out_r_39__N_1083[1] (\spi_data_out_r_39__N_1083[1] ), 
            .\spi_data_out_r_39__N_1083[26] (\spi_data_out_r_39__N_1083[26] ), 
            .spi_data_out_r_39__N_1398(spi_data_out_r_39__N_1398), .\spi_data_out_r_39__N_1083[25] (\spi_data_out_r_39__N_1083[25] ), 
            .\spi_data_out_r_39__N_1083[30] (\spi_data_out_r_39__N_1083[30] ), 
            .n30013(n30013), .\spi_data_out_r_39__N_2023[3] (\spi_data_out_r_39__N_2023[3] ), 
            .\SLO_buf[5]_adj_319 (\SLO_buf[5]_adj_642 ), .\spi_data_out_r_39__N_4419[1] (\spi_data_out_r_39__N_4419[1] ), 
            .\spi_data_out_r_39__N_2023[2] (\spi_data_out_r_39__N_2023[2] ), 
            .\spi_data_out_r_39__N_2023[1] (\spi_data_out_r_39__N_2023[1] ), 
            .\spi_data_out_r_39__N_1083[10] (\spi_data_out_r_39__N_1083[10] ), 
            .\spi_data_out_r_39__N_2023[0] (\spi_data_out_r_39__N_2023[0] ), 
            .\spi_data_out_r_39__N_2023[22] (\spi_data_out_r_39__N_2023[22] ), 
            .n30007(n30007), .n30016(n30016), .clk_enable_38(clk_enable_38), 
            .\spi_data_out_r_39__N_2023[21] (\spi_data_out_r_39__N_2023[21] ), 
            .n30020(n30020), .\spi_data_out_r_39__N_2023[31] (\spi_data_out_r_39__N_2023[31] ), 
            .clk_enable_227(clk_enable_227), .\spi_data_out_r_39__N_2023[30] (\spi_data_out_r_39__N_2023[30] ), 
            .\spi_data_out_r_39__N_2023[29] (\spi_data_out_r_39__N_2023[29] ), 
            .\spi_data_out_r_39__N_1083[28] (\spi_data_out_r_39__N_1083[28] ), 
            .\spi_data_out_r_39__N_2023[28] (\spi_data_out_r_39__N_2023[28] ), 
            .\spi_data_out_r_39__N_2023[27] (\spi_data_out_r_39__N_2023[27] ), 
            .\spi_data_out_r_39__N_1083[21] (\spi_data_out_r_39__N_1083[21] ), 
            .n22554(n22554), .pwm(pwm), .n4_adj_320(n4_adj_643), .\status_cntr[11] (\status_cntr[11] ), 
            .\spi_data_out_r_39__N_1083[0] (\spi_data_out_r_39__N_1083[0] ), 
            .spi_data_valid(spi_data_valid), .spi_data_out_r_39__N_2103(spi_data_out_r_39__N_2103), 
            .spi_data_out_r_39__N_1163(spi_data_out_r_39__N_1163), .\spi_data_out_r_39__N_2493[0] (\spi_data_out_r_39__N_2493[0] ), 
            .\spi_data_out_r_39__N_2493[31] (\spi_data_out_r_39__N_2493[31] ), 
            .\spi_data_out_r_39__N_2493[30] (\spi_data_out_r_39__N_2493[30] ), 
            .spi_data_out_r_39__N_1633(spi_data_out_r_39__N_1633), .spi_data_out_r_39__N_2573(spi_data_out_r_39__N_2573)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/spi_slave_top.v(203[4] 225[21])
    
endmodule
//
// Verilog Description of module wb_ctrl
//

module wb_ctrl (wb_cyc_i, clk, clk_enable_172, \wb_adr_i[0] , \address[0] , 
            wb_we_i, wb_we_i_N_344, wb_dat_i, wr_data, wb_sm, spi_cmd_start, 
            \address_7__N_549[1] , \address_7__N_565[1] , wr_en, wr_en_N_355, 
            \wb_adr_i[1] , \address[1] , \wb_adr_i[6] , n31069, rd_en, 
            n29) /* synthesis syn_module_defined=1 */ ;
    output wb_cyc_i;
    input clk;
    input clk_enable_172;
    output \wb_adr_i[0] ;
    input \address[0] ;
    output wb_we_i;
    input wb_we_i_N_344;
    output [7:0]wb_dat_i;
    input [7:0]wr_data;
    output wb_sm;
    input spi_cmd_start;
    input \address_7__N_549[1] ;
    output \address_7__N_565[1] ;
    input wr_en;
    output wr_en_N_355;
    output \wb_adr_i[1] ;
    input \address[1] ;
    output \wb_adr_i[6] ;
    input n31069;
    input rd_en;
    output n29;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    
    wire clk_enable_844, n11837, n30170;
    
    FD1P3AX wb_cyc_i_36 (.D(clk_enable_844), .SP(clk_enable_172), .CK(clk), 
            .Q(wb_cyc_i)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_cyc_i_36.GSR = "ENABLED";
    FD1P3AX wb_adr_i_i0 (.D(\address[0] ), .SP(clk_enable_844), .CK(clk), 
            .Q(\wb_adr_i[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_adr_i_i0.GSR = "ENABLED";
    FD1P3AX wb_we_i_38 (.D(wb_we_i_N_344), .SP(clk_enable_172), .CK(clk), 
            .Q(wb_we_i)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_we_i_38.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i0 (.D(wr_data[0]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i0.GSR = "ENABLED";
    FD1S3AX wb_sm_35 (.D(n11837), .CK(clk), .Q(wb_sm)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(83[11] 90[18])
    defparam wb_sm_35.GSR = "ENABLED";
    LUT4 i23561_4_lut (.A(spi_cmd_start), .B(n30170), .C(\address_7__N_549[1] ), 
         .D(wb_sm), .Z(\address_7__N_565[1] )) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(16[45:52])
    defparam i23561_4_lut.init = 16'ha022;
    LUT4 wr_en_I_0_1_lut (.A(wr_en), .Z(wr_en_N_355)) /* synthesis lut_function=(!(A)) */ ;   // c:/s_links/sources/wb_ctrl.v(129[44:50])
    defparam wr_en_I_0_1_lut.init = 16'h5555;
    FD1P3AX wb_adr_i_i1 (.D(\address[1] ), .SP(clk_enable_844), .CK(clk), 
            .Q(\wb_adr_i[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_adr_i_i1.GSR = "ENABLED";
    FD1P3AX wb_adr_i_i6 (.D(n31069), .SP(clk_enable_844), .CK(clk), .Q(\wb_adr_i[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_adr_i_i6.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i1 (.D(wr_data[1]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i1.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i2 (.D(wr_data[2]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i2.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i3 (.D(wr_data[3]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i3.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i4 (.D(wr_data[4]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i4.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i5 (.D(wr_data[5]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i5.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i6 (.D(wr_data[6]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i6.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i7 (.D(wr_data[7]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i7.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_770 (.A(wr_en), .B(rd_en), .Z(n30170)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_slave_top.v(53[44:49])
    defparam i1_2_lut_rep_770.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(wr_en), .B(rd_en), .C(wb_sm), 
         .D(\address_7__N_549[1] ), .Z(n11837)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // c:/s_links/sources/spi_slave_top.v(53[44:49])
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'h0efe;
    LUT4 i1_2_lut_rep_661_3_lut (.A(wr_en), .B(rd_en), .C(wb_sm), .Z(clk_enable_844)) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(53[44:49])
    defparam i1_2_lut_rep_661_3_lut.init = 16'h0e0e;
    LUT4 i61_3_lut_4_lut (.A(wr_en), .B(rd_en), .C(wb_sm), .D(\address_7__N_549[1] ), 
         .Z(n29)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // c:/s_links/sources/spi_slave_top.v(53[44:49])
    defparam i61_3_lut_4_lut.init = 16'hf101;
    
endmodule
//
// Verilog Description of module spi_slave_efb
//

module spi_slave_efb (clk, n30185, wb_cyc_i, wb_we_i, GND_net, \wb_adr_i[6] , 
            \wb_adr_i[1] , \wb_adr_i[0] , wb_dat_i, spi_scsn_c, wb_dat_o, 
            \address_7__N_549[1] , spi_mosi_oe, spi_mosi_o, spi_miso_oe, 
            spi_miso_o, spi_clk_oe, spi_clk_o, spi_mosi_i, spi_miso_i, 
            spi_clk_i, VCC_net, wb_sm, clk_enable_172) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input clk;
    input n30185;
    input wb_cyc_i;
    input wb_we_i;
    input GND_net;
    input \wb_adr_i[6] ;
    input \wb_adr_i[1] ;
    input \wb_adr_i[0] ;
    input [7:0]wb_dat_i;
    input spi_scsn_c;
    output [7:0]wb_dat_o;
    output \address_7__N_549[1] ;
    output spi_mosi_oe;
    output spi_mosi_o;
    output spi_miso_oe;
    output spi_miso_o;
    output spi_clk_oe;
    output spi_clk_o;
    input spi_mosi_i;
    input spi_miso_i;
    input spi_clk_i;
    input VCC_net;
    input wb_sm;
    output clk_enable_172;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire spi_clk_i /* synthesis is_clock=1 */ ;   // c:/s_links/sources/config_hex/ip/spi_slave_efb.v(34[10:19])
    
    EFB EFBInst_0 (.WBCLKI(clk), .WBRSTI(n30185), .WBCYCI(wb_cyc_i), .WBSTBI(wb_cyc_i), 
        .WBWEI(wb_we_i), .WBADRI0(\wb_adr_i[0] ), .WBADRI1(\wb_adr_i[1] ), 
        .WBADRI2(GND_net), .WBADRI3(\wb_adr_i[6] ), .WBADRI4(\wb_adr_i[6] ), 
        .WBADRI5(GND_net), .WBADRI6(\wb_adr_i[6] ), .WBADRI7(GND_net), 
        .WBDATI0(wb_dat_i[0]), .WBDATI1(wb_dat_i[1]), .WBDATI2(wb_dat_i[2]), 
        .WBDATI3(wb_dat_i[3]), .WBDATI4(wb_dat_i[4]), .WBDATI5(wb_dat_i[5]), 
        .WBDATI6(wb_dat_i[6]), .WBDATI7(wb_dat_i[7]), .I2C1SCLI(GND_net), 
        .I2C1SDAI(GND_net), .I2C2SCLI(GND_net), .I2C2SDAI(GND_net), .SPISCKI(spi_clk_i), 
        .SPIMISOI(spi_miso_i), .SPIMOSII(spi_mosi_i), .SPISCSN(spi_scsn_c), 
        .TCCLKI(GND_net), .TCRSTN(GND_net), .TCIC(GND_net), .UFMSN(VCC_net), 
        .PLL0DATI0(GND_net), .PLL0DATI1(GND_net), .PLL0DATI2(GND_net), 
        .PLL0DATI3(GND_net), .PLL0DATI4(GND_net), .PLL0DATI5(GND_net), 
        .PLL0DATI6(GND_net), .PLL0DATI7(GND_net), .PLL0ACKI(GND_net), 
        .PLL1DATI0(GND_net), .PLL1DATI1(GND_net), .PLL1DATI2(GND_net), 
        .PLL1DATI3(GND_net), .PLL1DATI4(GND_net), .PLL1DATI5(GND_net), 
        .PLL1DATI6(GND_net), .PLL1DATI7(GND_net), .PLL1ACKI(GND_net), 
        .WBDATO0(wb_dat_o[0]), .WBDATO1(wb_dat_o[1]), .WBDATO2(wb_dat_o[2]), 
        .WBDATO3(wb_dat_o[3]), .WBDATO4(wb_dat_o[4]), .WBDATO5(wb_dat_o[5]), 
        .WBDATO6(wb_dat_o[6]), .WBDATO7(wb_dat_o[7]), .WBACKO(\address_7__N_549[1] ), 
        .SPISCKO(spi_clk_o), .SPISCKEN(spi_clk_oe), .SPIMISOO(spi_miso_o), 
        .SPIMISOEN(spi_miso_oe), .SPIMOSIO(spi_mosi_o), .SPIMOSIEN(spi_mosi_oe)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=15, LSE_LLINE=162, LSE_RLINE=176 */ ;   // c:/s_links/sources/spi_slave_top.v(162[18] 176[15])
    defparam EFBInst_0.EFB_I2C1 = "DISABLED";
    defparam EFBInst_0.EFB_I2C2 = "DISABLED";
    defparam EFBInst_0.EFB_SPI = "ENABLED";
    defparam EFBInst_0.EFB_TC = "DISABLED";
    defparam EFBInst_0.EFB_TC_PORTMODE = "WB";
    defparam EFBInst_0.EFB_UFM = "DISABLED";
    defparam EFBInst_0.EFB_WB_CLK_FREQ = "100.0";
    defparam EFBInst_0.DEV_DENSITY = "4000L";
    defparam EFBInst_0.UFM_INIT_PAGES = 0;
    defparam EFBInst_0.UFM_INIT_START_PAGE = 0;
    defparam EFBInst_0.UFM_INIT_ALL_ZEROS = "ENABLED";
    defparam EFBInst_0.UFM_INIT_FILE_NAME = "NONE";
    defparam EFBInst_0.UFM_INIT_FILE_FORMAT = "HEX";
    defparam EFBInst_0.I2C1_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C2_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C1_SLAVE_ADDR = "0b1000001";
    defparam EFBInst_0.I2C2_SLAVE_ADDR = "0b1000010";
    defparam EFBInst_0.I2C1_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C2_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C1_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C2_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C1_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C2_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C1_WAKEUP = "DISABLED";
    defparam EFBInst_0.I2C2_WAKEUP = "DISABLED";
    defparam EFBInst_0.SPI_MODE = "SLAVE";
    defparam EFBInst_0.SPI_CLK_DIVIDER = 2;
    defparam EFBInst_0.SPI_LSB_FIRST = "DISABLED";
    defparam EFBInst_0.SPI_CLK_INV = "DISABLED";
    defparam EFBInst_0.SPI_PHASE_ADJ = "DISABLED";
    defparam EFBInst_0.SPI_SLAVE_HANDSHAKE = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXOVR = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXOVR = "DISABLED";
    defparam EFBInst_0.SPI_WAKEUP = "DISABLED";
    defparam EFBInst_0.TC_MODE = "CTCM";
    defparam EFBInst_0.TC_SCLK_SEL = "PCLOCK";
    defparam EFBInst_0.TC_CCLK_SEL = 1;
    defparam EFBInst_0.GSR = "ENABLED";
    defparam EFBInst_0.TC_TOP_SET = 65535;
    defparam EFBInst_0.TC_OCR_SET = 32767;
    defparam EFBInst_0.TC_OC_MODE = "TOGGLE";
    defparam EFBInst_0.TC_RESETN = "ENABLED";
    defparam EFBInst_0.TC_TOP_SEL = "OFF";
    defparam EFBInst_0.TC_OV_INT = "OFF";
    defparam EFBInst_0.TC_OCR_INT = "OFF";
    defparam EFBInst_0.TC_ICR_INT = "OFF";
    defparam EFBInst_0.TC_OVERFLOW = "DISABLED";
    defparam EFBInst_0.TC_ICAPTURE = "DISABLED";
    LUT4 i24014_2_lut_rep_737 (.A(\address_7__N_549[1] ), .B(wb_sm), .Z(clk_enable_172)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/spi_slave_top.v(162[18] 176[15])
    defparam i24014_2_lut_rep_737.init = 16'hbbbb;
    
endmodule
//
// Verilog Description of module spi_ctrl
//

module spi_ctrl (quad_buffer, quad_count, \spi_data_out_r_39__N_1083[31] , 
            spi_addr, spi_cmd, clk, \spi_data[0] , wb_dat_o, \spi_data_out_r_39__N_1083[29] , 
            wr_en_N_355, wr_data, \address[0] , rd_en, wr_en, spi_scsn_c, 
            \address_7__N_549[1] , \spi_data_out_r_39__N_1083[19] , \spi_data_out_r_39__N_1083[18] , 
            quad_buffer_adj_321, quad_count_adj_322, \spi_data_out_r_39__N_2023[26] , 
            n30198, n32, clear_intrpt_N_2717, \address_7__N_565[1] , 
            resetn_c, spi_addr_valid, n47, clear_intrpt_N_2930, clear_intrpt_N_2788, 
            clear_intrpt_N_2859, n47_adj_74, quad_buffer_adj_323, quad_count_adj_324, 
            \spi_data_out_r_39__N_2493[29] , \spi_data_out_r_39__N_2493[28] , 
            \spi_data_out_r_39__N_2493[27] , \spi_data_out_r_39__N_2493[26] , 
            n29997, n29991, \spi_data_out_r_39__N_2493[25] , \spi_data_out_r_39__N_2493[24] , 
            \spi_data_out_r_39__N_2493[23] , \spi_data_out_r_39__N_2493[22] , 
            \spi_data_out_r_39__N_2493[21] , \spi_data_out_r_39__N_2493[20] , 
            \spi_data_out_r_39__N_2493[19] , \spi_data[31] , \spi_data_out_r_39__N_2493[18] , 
            \spi_data_out_r_39__N_2493[17] , \spi_data_out_r_39__N_2493[16] , 
            \spi_data_out_r_39__N_2493[15] , \spi_data_out_r_39__N_2493[14] , 
            \spi_data_out_r_39__N_2493[13] , \spi_data_out_r_39__N_2493[12] , 
            \spi_data_out_r_39__N_2493[11] , \spi_data_out_r_39__N_2493[10] , 
            \spi_data[30] , \spi_data[29] , \spi_data[28] , \spi_data[27] , 
            \spi_data[26] , \spi_data[25] , \spi_data[24] , \spi_data[23] , 
            \spi_data[22] , \spi_data_out_r_39__N_2493[9] , \spi_data_out_r_39__N_2493[8] , 
            \spi_data[21] , \spi_data[20] , \spi_data[19] , \spi_data[18] , 
            \spi_data[17] , \spi_data_out_r_39__N_2493[7] , \spi_data[16] , 
            \spi_data[15] , \spi_data[14] , \spi_data[13] , \spi_data[12] , 
            \spi_data[11] , \spi_data[10] , \spi_data[9] , \spi_data[8] , 
            \spi_data[7] , \spi_data[6] , \spi_data[5] , \spi_data[4] , 
            \spi_data[3] , \spi_data_out_r_39__N_1083[9] , \spi_data[2] , 
            \spi_data[1] , \spi_data_out_r_39__N_1083[8] , \spi_data_out_r_39__N_2493[6] , 
            \spi_data_out_r_39__N_2493[5] , \spi_data_out_r_39__N_2493[4] , 
            \spi_data_out_r_39__N_2493[3] , \spi_data_out_r_39__N_2493[2] , 
            \spi_data_out_r_39__N_2493[1] , \spi_data_out_r_39__N_2023[20] , 
            quad_buffer_adj_325, quad_count_adj_326, \spi_data_out_r_39__N_2258[0] , 
            \spi_data_out_r_39__N_2258[31] , \spi_data_out_r_39__N_2258[30] , 
            \spi_data_out_r_39__N_2258[29] , \spi_data_out_r_39__N_2258[28] , 
            \spi_data_out_r_39__N_2258[27] , \spi_data_out_r_39__N_2258[26] , 
            n26779, \spi_data_out_r_39__N_2258[25] , \spi_data_out_r_39__N_2258[24] , 
            \spi_data_out_r_39__N_1083[22] , \spi_data_out_r_39__N_2258[23] , 
            \spi_data_out_r_39__N_2258[22] , \spi_data_out_r_39__N_2258[21] , 
            \spi_data_out_r_39__N_2258[20] , \spi_data_out_r_39__N_2258[19] , 
            \spi_data_out_r_39__N_2258[18] , n47_adj_203, \spi_data_out_r_39__N_2258[17] , 
            \spi_data_out_r_39__N_2258[16] , \spi_data_out_r_39__N_2258[15] , 
            \spi_data_out_r_39__N_2258[14] , \spi_data_out_r_39__N_2258[13] , 
            \spi_data_out_r_39__N_2258[12] , \spi_data_out_r_39__N_2258[11] , 
            \spi_data_out_r_39__N_2258[10] , \spi_data_out_r_39__N_2258[9] , 
            n30019, n47_adj_204, \spi_data_out_r_39__N_2258[8] , \address[1] , 
            \spi_data_out_r_39__N_2258[7] , n30027, n47_adj_205, \spi_data_out_r_39__N_2258[6] , 
            \spi_data_out_r_39__N_2258[5] , \spi_data_out_r_39__N_2258[4] , 
            \spi_data_out_r_39__N_2258[3] , \spi_data_out_r_39__N_1083[17] , 
            \spi_data_out_r_39__N_2258[2] , \spi_data_out_r_39__N_2023[19] , 
            \spi_data_out_r_39__N_2258[1] , \SLO_buf[4] , \SLO_buf[14] , 
            \spi_data_out_r_39__N_5105[0] , \SLO_buf[3] , \SLO_buf[9] , 
            \spi_data_out_r_39__N_5105[35] , \SLO_buf[2] , \SLO_buf[8] , 
            \spi_data_out_r_39__N_5105[34] , \SLO_buf[1] , \SLO_buf[7] , 
            \spi_data_out_r_39__N_5105[33] , quad_buffer_adj_327, quad_count_adj_328, 
            \spi_data_out_r_39__N_1553[0] , \spi_data_out_r_39__N_1553[31] , 
            \SLO_buf[0] , \SLO_buf[6] , \spi_data_out_r_39__N_5105[32] , 
            \SLO_buf[19] , \SLO_buf[29] , \spi_data_out_r_39__N_5105[15] , 
            \spi_data_out_r_39__N_1553[30] , \spi_data_out_r_39__N_1553[29] , 
            \spi_data_out_r_39__N_1553[28] , \spi_data_out_r_39__N_1553[27] , 
            \SLO_buf[18] , \SLO_buf[28] , \spi_data_out_r_39__N_5105[14] , 
            \spi_data_out_r_39__N_1553[26] , \SLO_buf[17] , \SLO_buf[27] , 
            \spi_data_out_r_39__N_5105[13] , \spi_data_out_r_39__N_2023[25] , 
            \spi_data_out_r_39__N_1553[25] , \spi_data_out_r_39__N_1553[24] , 
            wb_sm, wb_we_i_N_344, \SLO_buf[16] , \SLO_buf[26] , \spi_data_out_r_39__N_5105[12] , 
            \spi_data_out_r_39__N_1553[23] , \SLO_buf[15] , \SLO_buf[25] , 
            \spi_data_out_r_39__N_5105[11] , \SLO_buf[24] , \spi_data_out_r_39__N_5105[10] , 
            \spi_data_out_r_39__N_1553[22] , \SLO_buf[13] , \SLO_buf[23] , 
            \spi_data_out_r_39__N_5105[9] , \spi_data_out_r_39__N_1553[21] , 
            \spi_data_out_r_39__N_1553[20] , \spi_data_out_r_39__N_1553[19] , 
            \spi_data_out_r_39__N_1553[18] , \spi_data_out_r_39__N_1553[17] , 
            \spi_data_out_r_39__N_1553[16] , \spi_data_out_r_39__N_1083[16] , 
            \spi_data_out_r_39__N_1553[15] , \spi_data_out_r_39__N_1553[14] , 
            \spi_data_out_r_39__N_1553[13] , \spi_data_out_r_39__N_1083[15] , 
            GND_net, \SLO_buf[12] , \SLO_buf[22] , \spi_data_out_r_39__N_5105[8] , 
            \spi_data_out_r_39__N_1553[12] , \SLO_buf[11] , \SLO_buf[21] , 
            \spi_data_out_r_39__N_5105[7] , \spi_data_out_r_39__N_1553[11] , 
            \SLO_buf[10] , \SLO_buf[20] , \spi_data_out_r_39__N_5105[6] , 
            \spi_data_out_r_39__N_5105[5] , \spi_data_out_r_39__N_1553[10] , 
            \spi_data_out_r_39__N_5105[4] , \spi_data_out_r_39__N_1553[9] , 
            \spi_data_out_r_39__N_1553[8] , \spi_data_out_r_39__N_1553[7] , 
            \spi_data_out_r_39__N_1553[6] , \spi_data_out_r_39__N_5105[3] , 
            \spi_data_out_r_39__N_1553[5] , \spi_data_out_r_39__N_1553[4] , 
            \spi_data_out_r_39__N_1553[3] , \spi_data_out_r_39__N_2023[18] , 
            \spi_data_out_r_39__N_1553[2] , \spi_data_out_r_39__N_1553[1] , 
            n47_adj_270, spi_cmd_start, \spi_data_out_r_39__N_5105[2] , 
            \SLO_buf[5] , \spi_data_out_r_39__N_5105[1] , n29, spi_data_out_r_39__N_2338, 
            n47_adj_271, \spi_data_out_r_39__N_1083[14] , \spi_data_out_r_39__N_1083[13] , 
            n30102, \SLO_buf[4]_adj_272 , \SLO_buf[14]_adj_273 , \spi_data_out_r_39__N_4419[0] , 
            mem_rdata, \SLO_buf[3]_adj_274 , \SLO_buf[9]_adj_275 , \spi_data_out_r_39__N_4419[35] , 
            spi_data_out_r_39__N_4505, \spi_data_out_r_39__N_2023[17] , 
            \spi_data_out_r_39__N_2023[16] , \spi_data_out_r_39__N_1083[7] , 
            \spi_data_out_r_39__N_1083[6] , \spi_data_out_r_39__N_1083[20] , 
            \spi_data_out_r_39__N_2023[15] , \status_cntr[12] , n25212, 
            \SLO_buf[2]_adj_276 , \SLO_buf[8]_adj_277 , \spi_data_out_r_39__N_4419[34] , 
            \spi_data_out_r_39__N_2023[14] , \SLO_buf[1]_adj_278 , \SLO_buf[7]_adj_279 , 
            \spi_data_out_r_39__N_4419[33] , \SLO_buf[0]_adj_280 , \SLO_buf[6]_adj_281 , 
            \spi_data_out_r_39__N_4419[32] , clear_intrpt_N_3072, \spi_data_out_r_39__N_2023[13] , 
            \SLO_buf[19]_adj_282 , \SLO_buf[29]_adj_283 , \spi_data_out_r_39__N_4419[15] , 
            \spi_data_out_r_39__N_1083[5] , \spi_data_out_r_39__N_1083[4] , 
            \spi_data_out_r_39__N_2023[12] , \SLO_buf[18]_adj_284 , \SLO_buf[28]_adj_285 , 
            \spi_data_out_r_39__N_4419[14] , \SLO_buf[17]_adj_286 , \SLO_buf[27]_adj_287 , 
            \spi_data_out_r_39__N_4419[13] , \spi_data_out_r_39__N_1083[12] , 
            spi_data_out_r_39__N_4848, \spi_data_out_r_39__N_1083[3] , \spi_data_out_r_39__N_1083[2] , 
            \spi_data_out_r_39__N_2023[11] , \SLO_buf[16]_adj_288 , \SLO_buf[26]_adj_289 , 
            \spi_data_out_r_39__N_4419[12] , \spi_data_out_r_39__N_2023[10] , 
            \SLO_buf[15]_adj_290 , \SLO_buf[25]_adj_291 , \spi_data_out_r_39__N_4419[11] , 
            \SLO_buf[24]_adj_292 , \spi_data_out_r_39__N_4419[10] , \SLO_buf[13]_adj_293 , 
            \SLO_buf[23]_adj_294 , \spi_data_out_r_39__N_4419[9] , \SLO_buf[12]_adj_295 , 
            \SLO_buf[22]_adj_296 , \spi_data_out_r_39__N_4419[8] , n30185, 
            n25885, n30087, \quad_homing[1] , n1, spi_sdo_valid, clk_enable_963, 
            n30010, \spi_addr_r[0] , clk_enable_686, spi_cmd_valid, 
            spi_scsn_dly, clk_enable_776, n26077, n24066, n30062, 
            clk_enable_260, clear_intrpt, intrpt_out_N_2642, clear_intrpt_adj_297, 
            intrpt_out_N_3068, n28540, n30035, n23537, clk_enable_263, 
            quad_set_valid_N_1158, clk_enable_807, n20598, n8400, n12467, 
            n20647, n18654, n12435, n4, n30070, n26873, clk_enable_320, 
            n25877, n30075, \quad_homing[1]_adj_298 , n1_adj_299, n30199, 
            n23916, n26821, clk_enable_684, n26089, n26091, clk_enable_255, 
            EM_STOP, clk_enable_259, n29996, clk_enable_23, n26947, 
            clk_enable_253, pwm_out_N_3169, pwm_out_N_3153, clk_enable_15, 
            \spi_addr_r[7] , n26107, n30214, n26113, clear_intrpt_adj_300, 
            intrpt_out_N_2997, n25993, clk_enable_687, n30045, n28524, 
            clk_enable_759, clk_enable_48, clk_enable_624, n30033, n23526, 
            clk_enable_727, n11008, pwm_out_1_N_6491, clk_enable_613, 
            spi_sdo_valid_N_296, clk_enable_961, n30011, n26957, clk_enable_520, 
            n28364, n24065, n26033, clk_enable_232, clk_enable_254, 
            n29995, clk_enable_28, n28514, n26563, clk_enable_226, 
            clk_enable_639, clk_enable_228, pwm_out_3_N_6530, clk_enable_1105, 
            pwm_out_4_N_6549, clk_enable_1107, n26841, n26843, clk_enable_757, 
            n26023, n28366, clk_enable_245, pwm_out_2_N_6511, clk_enable_22, 
            n30022, n26415, clk_enable_488, n26633, clk_enable_641, 
            n25833, clk_enable_638, n30036, n26435, clk_enable_959, 
            n18440, n26249, clk_enable_235, clear_intrpt_adj_301, intrpt_out_N_2713, 
            n57, reset_r_N_4129, clk_enable_761, n30080, n29998, n26539, 
            clk_enable_738, n25881, n30095, \quad_homing[1]_adj_302 , 
            n1_adj_303, n28516, n26515, clk_enable_652, quad_set_valid_N_2098, 
            clk_enable_683, clk_enable_211, n2109, n25893, n30055, 
            \quad_homing[1]_adj_304 , n1_adj_305, n25869, n30043, \quad_homing[1]_adj_306 , 
            n1_adj_307, n25873, n30091, \quad_homing[1]_adj_308 , n1_adj_309, 
            n28476, n26059, clk_enable_32, clear_intrpt_adj_310, intrpt_out_N_2855, 
            clk_enable_178, clear_intrpt_adj_311, intrpt_out_N_2784, quad_set_valid_N_1393, 
            clk_enable_842, n27013, clk_enable_627, n26233, clk_enable_234, 
            quad_set_valid_N_2333, clk_enable_315, \SLO_buf[11]_adj_312 , 
            \SLO_buf[21]_adj_313 , \spi_data_out_r_39__N_4419[7] , clk_enable_256, 
            n29999, clk_enable_12, n26587, clk_enable_749, clk_enable_388, 
            n26207, clk_enable_898, clk_enable_180, n18, n2193, \SLO_buf[10]_adj_314 , 
            \SLO_buf[20]_adj_315 , \spi_data_out_r_39__N_4419[6] , clk_enable_244, 
            clear_intrpt_adj_316, intrpt_out_N_2926, pwm_out_1_N_6306, 
            clk_100k_enable_1, n25889, n30083, \quad_homing[1]_adj_317 , 
            n1_adj_318, clk_enable_595, n30039, \spi_data_out_r_39__N_2023[9] , 
            \spi_data_out_r_39__N_1083[24] , clear_intrpt_N_3001, \spi_data_out_r_39__N_2023[8] , 
            \spi_data_out_r_39__N_1083[11] , \spi_data_out_r_39__N_2023[7] , 
            \spi_data_out_r_39__N_1083[27] , \spi_data_out_r_39__N_4419[5] , 
            \spi_data_out_r_39__N_4419[4] , \spi_data_out_r_39__N_2023[6] , 
            n27095, spi_data_out_r_39__N_1868, n29992, \spi_data_out_r_39__N_4419[3] , 
            \spi_data_out_r_39__N_2023[5] , \spi_data_out_r_39__N_2023[24] , 
            \spi_data_out_r_39__N_4419[2] , n28452, spi_data_out_r_39__N_5191, 
            spi_data_out_r_39__N_5534, spi_data_out_r_39__N_5877, \spi_data_out_r_39__N_1083[23] , 
            spi_data_out_r_39__N_6220, \spi_data_out_r_39__N_2023[4] , \spi_data_out_r_39__N_2023[23] , 
            \spi_data_out_r_39__N_1083[1] , \spi_data_out_r_39__N_1083[26] , 
            spi_data_out_r_39__N_1398, \spi_data_out_r_39__N_1083[25] , 
            \spi_data_out_r_39__N_1083[30] , n30013, \spi_data_out_r_39__N_2023[3] , 
            \SLO_buf[5]_adj_319 , \spi_data_out_r_39__N_4419[1] , \spi_data_out_r_39__N_2023[2] , 
            \spi_data_out_r_39__N_2023[1] , \spi_data_out_r_39__N_1083[10] , 
            \spi_data_out_r_39__N_2023[0] , \spi_data_out_r_39__N_2023[22] , 
            n30007, n30016, clk_enable_38, \spi_data_out_r_39__N_2023[21] , 
            n30020, \spi_data_out_r_39__N_2023[31] , clk_enable_227, \spi_data_out_r_39__N_2023[30] , 
            \spi_data_out_r_39__N_2023[29] , \spi_data_out_r_39__N_1083[28] , 
            \spi_data_out_r_39__N_2023[28] , \spi_data_out_r_39__N_2023[27] , 
            \spi_data_out_r_39__N_1083[21] , n22554, pwm, n4_adj_320, 
            \status_cntr[11] , \spi_data_out_r_39__N_1083[0] , spi_data_valid, 
            spi_data_out_r_39__N_2103, spi_data_out_r_39__N_1163, \spi_data_out_r_39__N_2493[0] , 
            \spi_data_out_r_39__N_2493[31] , \spi_data_out_r_39__N_2493[30] , 
            spi_data_out_r_39__N_1633, spi_data_out_r_39__N_2573) /* synthesis syn_module_defined=1 */ ;
    input [31:0]quad_buffer;
    input [31:0]quad_count;
    output \spi_data_out_r_39__N_1083[31] ;
    output [7:0]spi_addr;
    output [15:0]spi_cmd;
    input clk;
    output \spi_data[0] ;
    input [7:0]wb_dat_o;
    output \spi_data_out_r_39__N_1083[29] ;
    input wr_en_N_355;
    output [7:0]wr_data;
    output \address[0] ;
    output rd_en;
    output wr_en;
    input spi_scsn_c;
    input \address_7__N_549[1] ;
    output \spi_data_out_r_39__N_1083[19] ;
    output \spi_data_out_r_39__N_1083[18] ;
    input [31:0]quad_buffer_adj_321;
    input [31:0]quad_count_adj_322;
    output \spi_data_out_r_39__N_2023[26] ;
    output n30198;
    output n32;
    output clear_intrpt_N_2717;
    input \address_7__N_565[1] ;
    input resetn_c;
    output spi_addr_valid;
    output n47;
    output clear_intrpt_N_2930;
    output clear_intrpt_N_2788;
    output clear_intrpt_N_2859;
    output n47_adj_74;
    input [31:0]quad_buffer_adj_323;
    input [31:0]quad_count_adj_324;
    output \spi_data_out_r_39__N_2493[29] ;
    output \spi_data_out_r_39__N_2493[28] ;
    output \spi_data_out_r_39__N_2493[27] ;
    output \spi_data_out_r_39__N_2493[26] ;
    output n29997;
    output n29991;
    output \spi_data_out_r_39__N_2493[25] ;
    output \spi_data_out_r_39__N_2493[24] ;
    output \spi_data_out_r_39__N_2493[23] ;
    output \spi_data_out_r_39__N_2493[22] ;
    output \spi_data_out_r_39__N_2493[21] ;
    output \spi_data_out_r_39__N_2493[20] ;
    output \spi_data_out_r_39__N_2493[19] ;
    output \spi_data[31] ;
    output \spi_data_out_r_39__N_2493[18] ;
    output \spi_data_out_r_39__N_2493[17] ;
    output \spi_data_out_r_39__N_2493[16] ;
    output \spi_data_out_r_39__N_2493[15] ;
    output \spi_data_out_r_39__N_2493[14] ;
    output \spi_data_out_r_39__N_2493[13] ;
    output \spi_data_out_r_39__N_2493[12] ;
    output \spi_data_out_r_39__N_2493[11] ;
    output \spi_data_out_r_39__N_2493[10] ;
    output \spi_data[30] ;
    output \spi_data[29] ;
    output \spi_data[28] ;
    output \spi_data[27] ;
    output \spi_data[26] ;
    output \spi_data[25] ;
    output \spi_data[24] ;
    output \spi_data[23] ;
    output \spi_data[22] ;
    output \spi_data_out_r_39__N_2493[9] ;
    output \spi_data_out_r_39__N_2493[8] ;
    output \spi_data[21] ;
    output \spi_data[20] ;
    output \spi_data[19] ;
    output \spi_data[18] ;
    output \spi_data[17] ;
    output \spi_data_out_r_39__N_2493[7] ;
    output \spi_data[16] ;
    output \spi_data[15] ;
    output \spi_data[14] ;
    output \spi_data[13] ;
    output \spi_data[12] ;
    output \spi_data[11] ;
    output \spi_data[10] ;
    output \spi_data[9] ;
    output \spi_data[8] ;
    output \spi_data[7] ;
    output \spi_data[6] ;
    output \spi_data[5] ;
    output \spi_data[4] ;
    output \spi_data[3] ;
    output \spi_data_out_r_39__N_1083[9] ;
    output \spi_data[2] ;
    output \spi_data[1] ;
    output \spi_data_out_r_39__N_1083[8] ;
    output \spi_data_out_r_39__N_2493[6] ;
    output \spi_data_out_r_39__N_2493[5] ;
    output \spi_data_out_r_39__N_2493[4] ;
    output \spi_data_out_r_39__N_2493[3] ;
    output \spi_data_out_r_39__N_2493[2] ;
    output \spi_data_out_r_39__N_2493[1] ;
    output \spi_data_out_r_39__N_2023[20] ;
    input [31:0]quad_buffer_adj_325;
    input [31:0]quad_count_adj_326;
    output \spi_data_out_r_39__N_2258[0] ;
    output \spi_data_out_r_39__N_2258[31] ;
    output \spi_data_out_r_39__N_2258[30] ;
    output \spi_data_out_r_39__N_2258[29] ;
    output \spi_data_out_r_39__N_2258[28] ;
    output \spi_data_out_r_39__N_2258[27] ;
    output \spi_data_out_r_39__N_2258[26] ;
    output n26779;
    output \spi_data_out_r_39__N_2258[25] ;
    output \spi_data_out_r_39__N_2258[24] ;
    output \spi_data_out_r_39__N_1083[22] ;
    output \spi_data_out_r_39__N_2258[23] ;
    output \spi_data_out_r_39__N_2258[22] ;
    output \spi_data_out_r_39__N_2258[21] ;
    output \spi_data_out_r_39__N_2258[20] ;
    output \spi_data_out_r_39__N_2258[19] ;
    output \spi_data_out_r_39__N_2258[18] ;
    output n47_adj_203;
    output \spi_data_out_r_39__N_2258[17] ;
    output \spi_data_out_r_39__N_2258[16] ;
    output \spi_data_out_r_39__N_2258[15] ;
    output \spi_data_out_r_39__N_2258[14] ;
    output \spi_data_out_r_39__N_2258[13] ;
    output \spi_data_out_r_39__N_2258[12] ;
    output \spi_data_out_r_39__N_2258[11] ;
    output \spi_data_out_r_39__N_2258[10] ;
    output \spi_data_out_r_39__N_2258[9] ;
    output n30019;
    output n47_adj_204;
    output \spi_data_out_r_39__N_2258[8] ;
    output \address[1] ;
    output \spi_data_out_r_39__N_2258[7] ;
    output n30027;
    output n47_adj_205;
    output \spi_data_out_r_39__N_2258[6] ;
    output \spi_data_out_r_39__N_2258[5] ;
    output \spi_data_out_r_39__N_2258[4] ;
    output \spi_data_out_r_39__N_2258[3] ;
    output \spi_data_out_r_39__N_1083[17] ;
    output \spi_data_out_r_39__N_2258[2] ;
    output \spi_data_out_r_39__N_2023[19] ;
    output \spi_data_out_r_39__N_2258[1] ;
    input \SLO_buf[4] ;
    input \SLO_buf[14] ;
    output \spi_data_out_r_39__N_5105[0] ;
    input \SLO_buf[3] ;
    input \SLO_buf[9] ;
    output \spi_data_out_r_39__N_5105[35] ;
    input \SLO_buf[2] ;
    input \SLO_buf[8] ;
    output \spi_data_out_r_39__N_5105[34] ;
    input \SLO_buf[1] ;
    input \SLO_buf[7] ;
    output \spi_data_out_r_39__N_5105[33] ;
    input [31:0]quad_buffer_adj_327;
    input [31:0]quad_count_adj_328;
    output \spi_data_out_r_39__N_1553[0] ;
    output \spi_data_out_r_39__N_1553[31] ;
    input \SLO_buf[0] ;
    input \SLO_buf[6] ;
    output \spi_data_out_r_39__N_5105[32] ;
    input \SLO_buf[19] ;
    input \SLO_buf[29] ;
    output \spi_data_out_r_39__N_5105[15] ;
    output \spi_data_out_r_39__N_1553[30] ;
    output \spi_data_out_r_39__N_1553[29] ;
    output \spi_data_out_r_39__N_1553[28] ;
    output \spi_data_out_r_39__N_1553[27] ;
    input \SLO_buf[18] ;
    input \SLO_buf[28] ;
    output \spi_data_out_r_39__N_5105[14] ;
    output \spi_data_out_r_39__N_1553[26] ;
    input \SLO_buf[17] ;
    input \SLO_buf[27] ;
    output \spi_data_out_r_39__N_5105[13] ;
    output \spi_data_out_r_39__N_2023[25] ;
    output \spi_data_out_r_39__N_1553[25] ;
    output \spi_data_out_r_39__N_1553[24] ;
    input wb_sm;
    output wb_we_i_N_344;
    input \SLO_buf[16] ;
    input \SLO_buf[26] ;
    output \spi_data_out_r_39__N_5105[12] ;
    output \spi_data_out_r_39__N_1553[23] ;
    input \SLO_buf[15] ;
    input \SLO_buf[25] ;
    output \spi_data_out_r_39__N_5105[11] ;
    input \SLO_buf[24] ;
    output \spi_data_out_r_39__N_5105[10] ;
    output \spi_data_out_r_39__N_1553[22] ;
    input \SLO_buf[13] ;
    input \SLO_buf[23] ;
    output \spi_data_out_r_39__N_5105[9] ;
    output \spi_data_out_r_39__N_1553[21] ;
    output \spi_data_out_r_39__N_1553[20] ;
    output \spi_data_out_r_39__N_1553[19] ;
    output \spi_data_out_r_39__N_1553[18] ;
    output \spi_data_out_r_39__N_1553[17] ;
    output \spi_data_out_r_39__N_1553[16] ;
    output \spi_data_out_r_39__N_1083[16] ;
    output \spi_data_out_r_39__N_1553[15] ;
    output \spi_data_out_r_39__N_1553[14] ;
    output \spi_data_out_r_39__N_1553[13] ;
    output \spi_data_out_r_39__N_1083[15] ;
    input GND_net;
    input \SLO_buf[12] ;
    input \SLO_buf[22] ;
    output \spi_data_out_r_39__N_5105[8] ;
    output \spi_data_out_r_39__N_1553[12] ;
    input \SLO_buf[11] ;
    input \SLO_buf[21] ;
    output \spi_data_out_r_39__N_5105[7] ;
    output \spi_data_out_r_39__N_1553[11] ;
    input \SLO_buf[10] ;
    input \SLO_buf[20] ;
    output \spi_data_out_r_39__N_5105[6] ;
    output \spi_data_out_r_39__N_5105[5] ;
    output \spi_data_out_r_39__N_1553[10] ;
    output \spi_data_out_r_39__N_5105[4] ;
    output \spi_data_out_r_39__N_1553[9] ;
    output \spi_data_out_r_39__N_1553[8] ;
    output \spi_data_out_r_39__N_1553[7] ;
    output \spi_data_out_r_39__N_1553[6] ;
    output \spi_data_out_r_39__N_5105[3] ;
    output \spi_data_out_r_39__N_1553[5] ;
    output \spi_data_out_r_39__N_1553[4] ;
    output \spi_data_out_r_39__N_1553[3] ;
    output \spi_data_out_r_39__N_2023[18] ;
    output \spi_data_out_r_39__N_1553[2] ;
    output \spi_data_out_r_39__N_1553[1] ;
    output n47_adj_270;
    output spi_cmd_start;
    output \spi_data_out_r_39__N_5105[2] ;
    input \SLO_buf[5] ;
    output \spi_data_out_r_39__N_5105[1] ;
    input n29;
    output spi_data_out_r_39__N_2338;
    output n47_adj_271;
    output \spi_data_out_r_39__N_1083[14] ;
    output \spi_data_out_r_39__N_1083[13] ;
    output n30102;
    input \SLO_buf[4]_adj_272 ;
    input \SLO_buf[14]_adj_273 ;
    output \spi_data_out_r_39__N_4419[0] ;
    input [7:0]mem_rdata;
    input \SLO_buf[3]_adj_274 ;
    input \SLO_buf[9]_adj_275 ;
    output \spi_data_out_r_39__N_4419[35] ;
    output spi_data_out_r_39__N_4505;
    output \spi_data_out_r_39__N_2023[17] ;
    output \spi_data_out_r_39__N_2023[16] ;
    output \spi_data_out_r_39__N_1083[7] ;
    output \spi_data_out_r_39__N_1083[6] ;
    output \spi_data_out_r_39__N_1083[20] ;
    output \spi_data_out_r_39__N_2023[15] ;
    input \status_cntr[12] ;
    output n25212;
    input \SLO_buf[2]_adj_276 ;
    input \SLO_buf[8]_adj_277 ;
    output \spi_data_out_r_39__N_4419[34] ;
    output \spi_data_out_r_39__N_2023[14] ;
    input \SLO_buf[1]_adj_278 ;
    input \SLO_buf[7]_adj_279 ;
    output \spi_data_out_r_39__N_4419[33] ;
    input \SLO_buf[0]_adj_280 ;
    input \SLO_buf[6]_adj_281 ;
    output \spi_data_out_r_39__N_4419[32] ;
    output clear_intrpt_N_3072;
    output \spi_data_out_r_39__N_2023[13] ;
    input \SLO_buf[19]_adj_282 ;
    input \SLO_buf[29]_adj_283 ;
    output \spi_data_out_r_39__N_4419[15] ;
    output \spi_data_out_r_39__N_1083[5] ;
    output \spi_data_out_r_39__N_1083[4] ;
    output \spi_data_out_r_39__N_2023[12] ;
    input \SLO_buf[18]_adj_284 ;
    input \SLO_buf[28]_adj_285 ;
    output \spi_data_out_r_39__N_4419[14] ;
    input \SLO_buf[17]_adj_286 ;
    input \SLO_buf[27]_adj_287 ;
    output \spi_data_out_r_39__N_4419[13] ;
    output \spi_data_out_r_39__N_1083[12] ;
    output spi_data_out_r_39__N_4848;
    output \spi_data_out_r_39__N_1083[3] ;
    output \spi_data_out_r_39__N_1083[2] ;
    output \spi_data_out_r_39__N_2023[11] ;
    input \SLO_buf[16]_adj_288 ;
    input \SLO_buf[26]_adj_289 ;
    output \spi_data_out_r_39__N_4419[12] ;
    output \spi_data_out_r_39__N_2023[10] ;
    input \SLO_buf[15]_adj_290 ;
    input \SLO_buf[25]_adj_291 ;
    output \spi_data_out_r_39__N_4419[11] ;
    input \SLO_buf[24]_adj_292 ;
    output \spi_data_out_r_39__N_4419[10] ;
    input \SLO_buf[13]_adj_293 ;
    input \SLO_buf[23]_adj_294 ;
    output \spi_data_out_r_39__N_4419[9] ;
    input \SLO_buf[12]_adj_295 ;
    input \SLO_buf[22]_adj_296 ;
    output \spi_data_out_r_39__N_4419[8] ;
    output n30185;
    input n25885;
    input n30087;
    input \quad_homing[1] ;
    output n1;
    input spi_sdo_valid;
    output clk_enable_963;
    input n30010;
    input \spi_addr_r[0] ;
    output clk_enable_686;
    output spi_cmd_valid;
    input spi_scsn_dly;
    output clk_enable_776;
    input n26077;
    input n24066;
    input n30062;
    output clk_enable_260;
    input clear_intrpt;
    output intrpt_out_N_2642;
    input clear_intrpt_adj_297;
    output intrpt_out_N_3068;
    input n28540;
    input n30035;
    input n23537;
    output clk_enable_263;
    input quad_set_valid_N_1158;
    output clk_enable_807;
    input n20598;
    output n8400;
    input n12467;
    input n20647;
    input n18654;
    output n12435;
    input n4;
    input n30070;
    input n26873;
    output clk_enable_320;
    input n25877;
    input n30075;
    input \quad_homing[1]_adj_298 ;
    output n1_adj_299;
    input n30199;
    input n23916;
    input n26821;
    output clk_enable_684;
    input n26089;
    input n26091;
    output clk_enable_255;
    input EM_STOP;
    input clk_enable_259;
    input n29996;
    output clk_enable_23;
    input n26947;
    output clk_enable_253;
    input pwm_out_N_3169;
    input pwm_out_N_3153;
    output clk_enable_15;
    input \spi_addr_r[7] ;
    input n26107;
    input n30214;
    output n26113;
    input clear_intrpt_adj_300;
    output intrpt_out_N_2997;
    input n25993;
    output clk_enable_687;
    input n30045;
    input n28524;
    output clk_enable_759;
    input clk_enable_48;
    output clk_enable_624;
    input n30033;
    input n23526;
    output clk_enable_727;
    input n11008;
    input pwm_out_1_N_6491;
    output clk_enable_613;
    input spi_sdo_valid_N_296;
    output clk_enable_961;
    input n30011;
    input n26957;
    output clk_enable_520;
    input n28364;
    input n24065;
    input n26033;
    output clk_enable_232;
    input clk_enable_254;
    input n29995;
    output clk_enable_28;
    input n28514;
    input n26563;
    output clk_enable_226;
    output clk_enable_639;
    output clk_enable_228;
    input pwm_out_3_N_6530;
    output clk_enable_1105;
    input pwm_out_4_N_6549;
    output clk_enable_1107;
    input n26841;
    input n26843;
    output clk_enable_757;
    input n26023;
    input n28366;
    output clk_enable_245;
    input pwm_out_2_N_6511;
    output clk_enable_22;
    input n30022;
    input n26415;
    output clk_enable_488;
    input n26633;
    output clk_enable_641;
    input n25833;
    output clk_enable_638;
    input n30036;
    input n26435;
    output clk_enable_959;
    input n18440;
    input n26249;
    output clk_enable_235;
    input clear_intrpt_adj_301;
    output intrpt_out_N_2713;
    output n57;
    input reset_r_N_4129;
    output clk_enable_761;
    output n30080;
    output n29998;
    input n26539;
    output clk_enable_738;
    input n25881;
    input n30095;
    input \quad_homing[1]_adj_302 ;
    output n1_adj_303;
    input n28516;
    input n26515;
    output clk_enable_652;
    input quad_set_valid_N_2098;
    output clk_enable_683;
    output clk_enable_211;
    output n2109;
    input n25893;
    input n30055;
    input \quad_homing[1]_adj_304 ;
    output n1_adj_305;
    input n25869;
    input n30043;
    input \quad_homing[1]_adj_306 ;
    output n1_adj_307;
    input n25873;
    input n30091;
    input \quad_homing[1]_adj_308 ;
    output n1_adj_309;
    input n28476;
    input n26059;
    output clk_enable_32;
    input clear_intrpt_adj_310;
    output intrpt_out_N_2855;
    output clk_enable_178;
    input clear_intrpt_adj_311;
    output intrpt_out_N_2784;
    input quad_set_valid_N_1393;
    output clk_enable_842;
    input n27013;
    output clk_enable_627;
    input n26233;
    output clk_enable_234;
    input quad_set_valid_N_2333;
    output clk_enable_315;
    input \SLO_buf[11]_adj_312 ;
    input \SLO_buf[21]_adj_313 ;
    output \spi_data_out_r_39__N_4419[7] ;
    input clk_enable_256;
    input n29999;
    output clk_enable_12;
    input n26587;
    output clk_enable_749;
    output clk_enable_388;
    input n26207;
    output clk_enable_898;
    output clk_enable_180;
    input n18;
    output n2193;
    input \SLO_buf[10]_adj_314 ;
    input \SLO_buf[20]_adj_315 ;
    output \spi_data_out_r_39__N_4419[6] ;
    output clk_enable_244;
    input clear_intrpt_adj_316;
    output intrpt_out_N_2926;
    input pwm_out_1_N_6306;
    output clk_100k_enable_1;
    input n25889;
    input n30083;
    input \quad_homing[1]_adj_317 ;
    output n1_adj_318;
    output clk_enable_595;
    output n30039;
    output \spi_data_out_r_39__N_2023[9] ;
    output \spi_data_out_r_39__N_1083[24] ;
    output clear_intrpt_N_3001;
    output \spi_data_out_r_39__N_2023[8] ;
    output \spi_data_out_r_39__N_1083[11] ;
    output \spi_data_out_r_39__N_2023[7] ;
    output \spi_data_out_r_39__N_1083[27] ;
    output \spi_data_out_r_39__N_4419[5] ;
    output \spi_data_out_r_39__N_4419[4] ;
    output \spi_data_out_r_39__N_2023[6] ;
    output n27095;
    output spi_data_out_r_39__N_1868;
    output n29992;
    output \spi_data_out_r_39__N_4419[3] ;
    output \spi_data_out_r_39__N_2023[5] ;
    output \spi_data_out_r_39__N_2023[24] ;
    output \spi_data_out_r_39__N_4419[2] ;
    output n28452;
    output spi_data_out_r_39__N_5191;
    output spi_data_out_r_39__N_5534;
    output spi_data_out_r_39__N_5877;
    output \spi_data_out_r_39__N_1083[23] ;
    output spi_data_out_r_39__N_6220;
    output \spi_data_out_r_39__N_2023[4] ;
    output \spi_data_out_r_39__N_2023[23] ;
    output \spi_data_out_r_39__N_1083[1] ;
    output \spi_data_out_r_39__N_1083[26] ;
    output spi_data_out_r_39__N_1398;
    output \spi_data_out_r_39__N_1083[25] ;
    output \spi_data_out_r_39__N_1083[30] ;
    output n30013;
    output \spi_data_out_r_39__N_2023[3] ;
    input \SLO_buf[5]_adj_319 ;
    output \spi_data_out_r_39__N_4419[1] ;
    output \spi_data_out_r_39__N_2023[2] ;
    output \spi_data_out_r_39__N_2023[1] ;
    output \spi_data_out_r_39__N_1083[10] ;
    output \spi_data_out_r_39__N_2023[0] ;
    output \spi_data_out_r_39__N_2023[22] ;
    input n30007;
    input n30016;
    output clk_enable_38;
    output \spi_data_out_r_39__N_2023[21] ;
    output n30020;
    output \spi_data_out_r_39__N_2023[31] ;
    output clk_enable_227;
    output \spi_data_out_r_39__N_2023[30] ;
    output \spi_data_out_r_39__N_2023[29] ;
    output \spi_data_out_r_39__N_1083[28] ;
    output \spi_data_out_r_39__N_2023[28] ;
    output \spi_data_out_r_39__N_2023[27] ;
    output \spi_data_out_r_39__N_1083[21] ;
    input n22554;
    input pwm;
    input n4_adj_320;
    input \status_cntr[11] ;
    output \spi_data_out_r_39__N_1083[0] ;
    output spi_data_valid;
    output spi_data_out_r_39__N_2103;
    output spi_data_out_r_39__N_1163;
    output \spi_data_out_r_39__N_2493[0] ;
    output \spi_data_out_r_39__N_2493[31] ;
    output \spi_data_out_r_39__N_2493[30] ;
    output spi_data_out_r_39__N_1633;
    output spi_data_out_r_39__N_2573;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    
    wire n23623, n30159, n27151;
    wire [3:0]spi_byte_cnt;   // c:/s_links/sources/spi_ctrl.v(74[13:25])
    
    wire clk_enable_915, n12446, n30182, clk_enable_584, n6196, mem_wr, 
        n11068, n30092, n30074, n28444, n30135, n26721, n23208, 
        n30212;
    wire [15:0]n1220;
    
    wire n26, n38, spi_cmd_start_reg_N_745, n22944;
    wire [7:0]n2;
    
    wire mem_rdata_update, n8127, clk_enable_756;
    wire [7:0]n672;
    
    wire spi_idle_N_747, spi_csn_buf0_p, spi_csn_buf2_p, spi_cmd_start_reg, 
        n30226, spi_idle, n12176;
    wire [7:0]address_7__N_359;
    
    wire rd_en_N_710, wr_en_N_697, spi_cmd_cnt, spi_cmd_cnt_N_749, n30221, 
        clk_enable_859, n30127, spi_data_valid_N_737, n30200, n27171, 
        n27169, n30169, n10255, n30017, n24822, n24802, n30217, 
        n11723, n28426, n26467, n26461, n30194, mem_rdata_update_N_729, 
        n8000, n11728;
    wire [1:0]n5327;
    
    wire n9392, n28577, n30223, n24505, spi_addr_valid_N_732, n7951, 
        n7957, n24758, n30123, n7963, n7965, n24465, spi_cmd_start_reg_N_746, 
        n7977, clk_enable_321, n26597, n26599, n30069, n30160, n26483, 
        n27215, n27197, n30084, n27157, n30101, n26445, n16817, 
        n29911, n29910, n29912, n27049, n30154, n27081, n32_adj_6711, 
        n28573, n30161, n16815, n24275, n30225, n27137, n30224, 
        clk_enable_561, clk_enable_569, clk_enable_577, n30157, n30158, 
        n30096, rd_en_N_717, n26715, n28290, n30147, n26771, n26641;
    wire [3:0]n21;
    
    wire n26655, n27065, n30145, n27057, n31067, n30173;
    wire [7:0]n37;
    
    wire n27037, n27027, n26355, n30026, n27077, n30156, n30136;
    wire [7:0]mem_burst_cnt;   // c:/s_links/sources/spi_ctrl.v(71[16:29])
    
    wire n23343, n18233, n27089, n27177, wr_en_N_701, n11758, clk_enable_867, 
        n28534, n25421, n12, n11759, n23860, n28508, n10254, n7970, 
        n24183, n6, n21900, n21899, n21898, n30193, n30093, n26653, 
        n21897, n23412, n24310, n23469, n26263, n30059, n30211, 
        n27127, n30197, n30216, n24198, n29985, n23360, n30054, 
        n27211, n30195, n21890;
    wire [7:0]n37_adj_7039;
    
    wire n21889, n21888, n21887, n12460, n30196, n27229, n27223, 
        clk_enable_1128, n27365, n30000, n28506, n25271, n27259, 
        n26013, n26015, n26007, n26011, n30222, n27143, n30012, 
        n27239, n27323, n27183, n27245, n1277, n26257, n24312, 
        n24466, n26661, n24197, n26765, n8019, n4382, n11727, 
        n26333, n30060, n25457, n26043, n8, n30113, clk_enable_1110, 
        n18232, clk_enable_1106, n18231;
    
    LUT4 mux_422_i32_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[31]), 
         .D(quad_count[31]), .Z(\spi_data_out_r_39__N_1083[31] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_4_lut (.A(spi_addr[0]), .B(spi_addr[1]), .C(spi_cmd[15]), 
         .D(spi_cmd[7]), .Z(n27151)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_3_lut_4_lut.init = 16'h0080;
    FD1P3IX spi_byte_cnt_1788__i0 (.D(n30182), .SP(clk_enable_915), .CD(n12446), 
            .CK(clk), .Q(spi_byte_cnt[0]));   // c:/s_links/sources/spi_ctrl.v(383[46:62])
    defparam spi_byte_cnt_1788__i0.GSR = "ENABLED";
    FD1P3IX spi_data__i0 (.D(wb_dat_o[0]), .SP(clk_enable_584), .CD(n6196), 
            .CK(clk), .Q(\spi_data[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i0.GSR = "ENABLED";
    FD1S3IX mem_wr_219 (.D(n30092), .CK(clk), .CD(n11068), .Q(mem_wr)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mem_wr_219.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut (.A(n30074), .B(n28444), .C(n30135), .D(n26721), 
         .Z(n23208)) /* synthesis lut_function=(!(A+!(B (C)+!B (C+(D))))) */ ;   // c:/s_links/sources/spi_ctrl.v(249[31] 252[34])
    defparam i1_4_lut_4_lut.init = 16'h5150;
    LUT4 i60_4_lut_4_lut (.A(n30074), .B(n30212), .C(n1220[10]), .D(n26), 
         .Z(n38)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/s_links/sources/spi_ctrl.v(249[31] 252[34])
    defparam i60_4_lut_4_lut.init = 16'h4f40;
    FD1S3AY main_sm_FSM_i1 (.D(n22944), .CK(clk), .Q(spi_cmd_start_reg_N_745));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i1.GSR = "ENABLED";
    FD1P3AX mem_addr_1792__i0 (.D(n2[0]), .SP(clk_enable_915), .CK(clk), 
            .Q(spi_addr[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_1792__i0.GSR = "ENABLED";
    LUT4 mux_422_i30_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[29]), 
         .D(quad_count[29]), .Z(\spi_data_out_r_39__N_1083[29] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i30_3_lut_4_lut.init = 16'hf1e0;
    FD1S3IX mem_rdata_update_206 (.D(n8127), .CK(clk), .CD(wr_en_N_355), 
            .Q(mem_rdata_update)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(79[9] 86[5])
    defparam mem_rdata_update_206.GSR = "DISABLED";
    FD1P3AX wr_data_i0_i0 (.D(n672[0]), .SP(clk_enable_756), .CK(clk), 
            .Q(wr_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i0.GSR = "ENABLED";
    FD1S3AY spi_csn_buf1_p_209 (.D(spi_csn_buf0_p), .CK(clk), .Q(spi_idle_N_747)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(103[11:44])
    defparam spi_csn_buf1_p_209.GSR = "ENABLED";
    FD1S3AY spi_csn_buf2_p_210 (.D(spi_idle_N_747), .CK(clk), .Q(spi_csn_buf2_p)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(110[11:44])
    defparam spi_csn_buf2_p_210.GSR = "ENABLED";
    FD1S3AX spi_cmd_start_reg_211 (.D(n30226), .CK(clk), .Q(spi_cmd_start_reg)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(117[11] 120[40])
    defparam spi_cmd_start_reg_211.GSR = "ENABLED";
    FD1S3AX spi_idle_212 (.D(n12176), .CK(clk), .Q(spi_idle)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(130[11] 133[31])
    defparam spi_idle_212.GSR = "ENABLED";
    FD1S3AY address_i1 (.D(address_7__N_359[0]), .CK(clk), .Q(\address[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam address_i1.GSR = "ENABLED";
    FD1S3AX rd_en_215 (.D(rd_en_N_710), .CK(clk), .Q(rd_en)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam rd_en_215.GSR = "ENABLED";
    FD1S3AX wr_en_216 (.D(wr_en_N_697), .CK(clk), .Q(wr_en)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_en_216.GSR = "ENABLED";
    FD1S3AX spi_cmd_cnt_228 (.D(spi_cmd_cnt_N_749), .CK(clk), .Q(spi_cmd_cnt)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_cnt_228.GSR = "ENABLED";
    FD1S3AY spi_csn_buf0_p_208 (.D(spi_scsn_c), .CK(clk), .Q(spi_csn_buf0_p)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(96[11:37])
    defparam spi_csn_buf0_p_208.GSR = "ENABLED";
    LUT4 i3740_4_lut_else_4_lut (.A(\address_7__N_549[1] ), .B(n1220[9]), 
         .C(wb_dat_o[3]), .Z(n30221)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i3740_4_lut_else_4_lut.init = 16'h8080;
    LUT4 mux_422_i20_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[19]), 
         .D(quad_count[19]), .Z(\spi_data_out_r_39__N_1083[19] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i20_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AY spi_cmd_i0_i0 (.D(wb_dat_o[0]), .SP(clk_enable_859), .CK(clk), 
            .Q(spi_cmd[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i0.GSR = "ENABLED";
    LUT4 mux_422_i19_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[18]), 
         .D(quad_count[18]), .Z(\spi_data_out_r_39__N_1083[18] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut (.A(spi_cmd[15]), .B(n30127), .C(spi_data_valid_N_737), 
         .Z(clk_enable_584)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_3_lut.init = 16'h4040;
    LUT4 mux_426_i27_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[26]), 
         .D(quad_count_adj_322[26]), .Z(\spi_data_out_r_39__N_2023[26] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut (.A(n27171), .B(n30198), .C(n32), .D(n27169), .Z(clear_intrpt_N_2717)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0200;
    LUT4 i2_2_lut_4_lut (.A(spi_idle), .B(n30169), .C(wb_dat_o[3]), .D(n1220[9]), 
         .Z(n10255)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:73])
    defparam i2_2_lut_4_lut.init = 16'hfe00;
    LUT4 i24017_2_lut_rep_617_4_lut (.A(spi_idle), .B(n30169), .C(wb_dat_o[3]), 
         .D(\address_7__N_549[1] ), .Z(n30017)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C (D))))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:73])
    defparam i24017_2_lut_rep_617_4_lut.init = 16'h01ff;
    LUT4 i1_4_lut_adj_593 (.A(spi_cmd_start_reg_N_745), .B(n30074), .C(\address_7__N_565[1] ), 
         .D(n24822), .Z(n22944)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_593.init = 16'hce0a;
    LUT4 i1_4_lut_adj_594 (.A(\address_7__N_549[1] ), .B(n11068), .C(n1220[5]), 
         .D(n24802), .Z(n24822)) /* synthesis lut_function=(A ((C+(D))+!B)+!A ((C)+!B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_594.init = 16'hfbf3;
    LUT4 i1_4_lut_adj_595 (.A(n1220[7]), .B(n30217), .C(n1220[11]), .D(n11723), 
         .Z(n24802)) /* synthesis lut_function=(A+(B (C)+!B (C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_595.init = 16'hfbfa;
    LUT4 i4_2_lut (.A(n1220[3]), .B(n1220[9]), .Z(n11723)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i23724_3_lut_4_lut (.A(n1220[4]), .B(n30135), .C(\address_7__N_549[1] ), 
         .D(n1220[10]), .Z(n28426)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i23724_3_lut_4_lut.init = 16'hefee;
    FD1P3AX mem_addr_1792__i7 (.D(n2[7]), .SP(clk_enable_915), .CK(clk), 
            .Q(spi_addr[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_1792__i7.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_596 (.A(n26467), .B(n30198), .C(n32), .D(n26461), 
         .Z(n23623)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_596.init = 16'hfffe;
    FD1P3AX mem_addr_1792__i6 (.D(n2[6]), .SP(clk_enable_915), .CK(clk), 
            .Q(spi_addr[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_1792__i6.GSR = "ENABLED";
    FD1P3AX mem_addr_1792__i5 (.D(n2[5]), .SP(clk_enable_915), .CK(clk), 
            .Q(spi_addr[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_1792__i5.GSR = "ENABLED";
    FD1P3AX mem_addr_1792__i4 (.D(n2[4]), .SP(clk_enable_915), .CK(clk), 
            .Q(spi_addr[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_1792__i4.GSR = "ENABLED";
    FD1P3AX mem_addr_1792__i3 (.D(n2[3]), .SP(clk_enable_915), .CK(clk), 
            .Q(spi_addr[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_1792__i3.GSR = "ENABLED";
    FD1P3AX mem_addr_1792__i2 (.D(n2[2]), .SP(clk_enable_915), .CK(clk), 
            .Q(spi_addr[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_1792__i2.GSR = "ENABLED";
    FD1P3AX mem_addr_1792__i1 (.D(n2[1]), .SP(clk_enable_915), .CK(clk), 
            .Q(spi_addr[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_1792__i1.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_597 (.A(n30194), .B(spi_cmd[2]), .C(spi_cmd[7]), 
         .D(spi_addr[1]), .Z(n26461)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_597.init = 16'hfffe;
    FD1S3AX main_sm_FSM_i13 (.D(n8000), .CK(clk), .Q(mem_rdata_update_N_729));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i13.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i12 (.D(n11728), .CK(clk), .Q(n1220[11]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i12.GSR = "ENABLED";
    PFUMX i5069 (.BLUT(n5327[1]), .ALUT(n9392), .C0(n28577), .Z(address_7__N_359[1]));
    FD1S3AX main_sm_FSM_i11 (.D(n30223), .CK(clk), .Q(n1220[10]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i11.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i10 (.D(n24505), .CK(clk), .Q(n1220[9]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i10.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i9 (.D(n7951), .CK(clk), .Q(spi_addr_valid_N_732));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i9.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i8 (.D(n7957), .CK(clk), .Q(n1220[7]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i8.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i7 (.D(n24758), .CK(clk), .Q(n1220[6]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i7.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i6 (.D(n30123), .CK(clk), .Q(n1220[5]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i6.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i5 (.D(n7963), .CK(clk), .Q(n1220[4]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i5.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i4 (.D(n7965), .CK(clk), .Q(n1220[3]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i4.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i3 (.D(n24465), .CK(clk), .Q(n1220[2]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i3.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i2 (.D(n7977), .CK(clk), .Q(spi_cmd_start_reg_N_746));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i2.GSR = "ENABLED";
    LUT4 i3803_2_lut (.A(mem_rdata_update_N_729), .B(resetn_c), .Z(n8127)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_ctrl.v(79[9] 86[5])
    defparam i3803_2_lut.init = 16'h8888;
    FD1P3AX spi_addr_valid_224 (.D(spi_addr_valid_N_732), .SP(clk_enable_321), 
            .CK(clk), .Q(spi_addr_valid)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_addr_valid_224.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_598 (.A(n26597), .B(n30198), .C(n26599), .D(n30069), 
         .Z(n47)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_598.init = 16'hfffe;
    LUT4 i1_2_lut (.A(spi_cmd[2]), .B(n32), .Z(n26597)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut.init = 16'hdddd;
    LUT4 i24126_2_lut_3_lut_4_lut (.A(spi_addr[1]), .B(n30160), .C(n26483), 
         .D(spi_cmd[2]), .Z(clear_intrpt_N_2930)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i24126_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_4_lut_adj_599 (.A(n27215), .B(n30198), .C(n27197), .D(n30084), 
         .Z(clear_intrpt_N_2788)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_4_lut_adj_599.init = 16'h0020;
    LUT4 i1_4_lut_adj_600 (.A(n27157), .B(n30198), .C(n32), .D(n30084), 
         .Z(clear_intrpt_N_2859)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_600.init = 16'h0002;
    LUT4 i1_4_lut_adj_601 (.A(n27151), .B(n30194), .C(n30101), .D(spi_cmd[2]), 
         .Z(n27157)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_601.init = 16'h0002;
    LUT4 i1_4_lut_adj_602 (.A(n26445), .B(n30198), .C(n26597), .D(spi_cmd[15]), 
         .Z(n16817)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_602.init = 16'hfeff;
    LUT4 i1_4_lut_adj_603 (.A(n30194), .B(n30084), .C(n30101), .D(spi_cmd[7]), 
         .Z(n26445)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_603.init = 16'hfffe;
    PFUMX i24369 (.BLUT(n29911), .ALUT(n29910), .C0(n30074), .Z(n29912));
    LUT4 i1_4_lut_adj_604 (.A(n27049), .B(n30198), .C(n30154), .D(n27081), 
         .Z(n47_adj_74)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_604.init = 16'hffef;
    PFUMX i57 (.BLUT(n38), .ALUT(n32_adj_6711), .C0(n28573), .Z(rd_en_N_710));
    LUT4 i1_4_lut_adj_605 (.A(n32), .B(n30194), .C(n30161), .D(n30160), 
         .Z(n27049)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_605.init = 16'hfffe;
    LUT4 mux_428_i30_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[29]), 
         .D(quad_count_adj_324[29]), .Z(\spi_data_out_r_39__N_2493[29] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i29_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[28]), 
         .D(quad_count_adj_324[28]), .Z(\spi_data_out_r_39__N_2493[28] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i28_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[27]), 
         .D(quad_count_adj_324[27]), .Z(\spi_data_out_r_39__N_2493[27] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i27_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[26]), 
         .D(quad_count_adj_324[26]), .Z(\spi_data_out_r_39__N_2493[26] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_rep_34_4_lut_4_lut_4_lut (.A(n29997), .B(spi_cmd[1]), .C(spi_addr[3]), 
         .D(spi_cmd[2]), .Z(n24275)) /* synthesis lut_function=(A+(B (C+(D))+!B (C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_rep_34_4_lut_4_lut_4_lut.init = 16'hfefb;
    LUT4 i1_2_lut_rep_591_3_lut (.A(spi_addr[0]), .B(spi_addr[1]), .C(n16817), 
         .Z(n29991)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_2_lut_rep_591_3_lut.init = 16'hf7f7;
    LUT4 i7817_4_lut_then_2_lut (.A(spi_idle_N_747), .B(spi_csn_buf2_p), 
         .Z(n30225)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/s_links/sources/spi_ctrl.v(117[11] 120[40])
    defparam i7817_4_lut_then_2_lut.init = 16'h4444;
    LUT4 mux_428_i26_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[25]), 
         .D(quad_count_adj_324[25]), .Z(\spi_data_out_r_39__N_2493[25] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i25_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[24]), 
         .D(quad_count_adj_324[24]), .Z(\spi_data_out_r_39__N_2493[24] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(spi_addr[0]), .B(spi_addr[1]), .C(spi_cmd[2]), 
         .D(spi_cmd[15]), .Z(n27137)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i7817_4_lut_else_2_lut (.A(spi_idle_N_747), .B(spi_csn_buf2_p), 
         .C(spi_cmd_start_reg_N_745), .D(spi_cmd_start_reg), .Z(n30224)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B+!(C+!(D))))) */ ;   // c:/s_links/sources/spi_ctrl.v(117[11] 120[40])
    defparam i7817_4_lut_else_2_lut.init = 16'h4d44;
    LUT4 mux_428_i24_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[23]), 
         .D(quad_count_adj_324[23]), .Z(\spi_data_out_r_39__N_2493[23] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i23_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[22]), 
         .D(quad_count_adj_324[22]), .Z(\spi_data_out_r_39__N_2493[22] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i22_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[21]), 
         .D(quad_count_adj_324[21]), .Z(\spi_data_out_r_39__N_2493[21] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i21_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[20]), 
         .D(quad_count_adj_324[20]), .Z(\spi_data_out_r_39__N_2493[20] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i20_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[19]), 
         .D(quad_count_adj_324[19]), .Z(\spi_data_out_r_39__N_2493[19] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i20_3_lut_4_lut.init = 16'hf1e0;
    FD1P3IX spi_data__i31 (.D(wb_dat_o[7]), .SP(clk_enable_561), .CD(n6196), 
            .CK(clk), .Q(\spi_data[31] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i31.GSR = "ENABLED";
    LUT4 mux_428_i19_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[18]), 
         .D(quad_count_adj_324[18]), .Z(\spi_data_out_r_39__N_2493[18] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i18_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[17]), 
         .D(quad_count_adj_324[17]), .Z(\spi_data_out_r_39__N_2493[17] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i17_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[16]), 
         .D(quad_count_adj_324[16]), .Z(\spi_data_out_r_39__N_2493[16] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i16_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[15]), 
         .D(quad_count_adj_324[15]), .Z(\spi_data_out_r_39__N_2493[15] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i15_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[14]), 
         .D(quad_count_adj_324[14]), .Z(\spi_data_out_r_39__N_2493[14] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i14_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[13]), 
         .D(quad_count_adj_324[13]), .Z(\spi_data_out_r_39__N_2493[13] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i13_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[12]), 
         .D(quad_count_adj_324[12]), .Z(\spi_data_out_r_39__N_2493[12] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i12_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[11]), 
         .D(quad_count_adj_324[11]), .Z(\spi_data_out_r_39__N_2493[11] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i11_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[10]), 
         .D(quad_count_adj_324[10]), .Z(\spi_data_out_r_39__N_2493[10] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i11_3_lut_4_lut.init = 16'hf1e0;
    FD1P3IX spi_data__i30 (.D(wb_dat_o[6]), .SP(clk_enable_561), .CD(n6196), 
            .CK(clk), .Q(\spi_data[30] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i30.GSR = "ENABLED";
    FD1P3IX spi_data__i29 (.D(wb_dat_o[5]), .SP(clk_enable_561), .CD(n6196), 
            .CK(clk), .Q(\spi_data[29] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i29.GSR = "ENABLED";
    FD1P3IX spi_data__i28 (.D(wb_dat_o[4]), .SP(clk_enable_561), .CD(n6196), 
            .CK(clk), .Q(\spi_data[28] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i28.GSR = "ENABLED";
    FD1P3IX spi_data__i27 (.D(wb_dat_o[3]), .SP(clk_enable_561), .CD(n6196), 
            .CK(clk), .Q(\spi_data[27] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i27.GSR = "ENABLED";
    FD1P3IX spi_data__i26 (.D(wb_dat_o[2]), .SP(clk_enable_561), .CD(n6196), 
            .CK(clk), .Q(\spi_data[26] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i26.GSR = "ENABLED";
    FD1P3IX spi_data__i25 (.D(wb_dat_o[1]), .SP(clk_enable_561), .CD(n6196), 
            .CK(clk), .Q(\spi_data[25] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i25.GSR = "ENABLED";
    FD1P3IX spi_data__i24 (.D(wb_dat_o[0]), .SP(clk_enable_561), .CD(n6196), 
            .CK(clk), .Q(\spi_data[24] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i24.GSR = "ENABLED";
    FD1P3IX spi_data__i23 (.D(wb_dat_o[7]), .SP(clk_enable_569), .CD(n6196), 
            .CK(clk), .Q(\spi_data[23] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i23.GSR = "ENABLED";
    FD1P3IX spi_data__i22 (.D(wb_dat_o[6]), .SP(clk_enable_569), .CD(n6196), 
            .CK(clk), .Q(\spi_data[22] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i22.GSR = "ENABLED";
    LUT4 mux_428_i10_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[9]), 
         .D(quad_count_adj_324[9]), .Z(\spi_data_out_r_39__N_2493[9] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i9_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[8]), 
         .D(quad_count_adj_324[8]), .Z(\spi_data_out_r_39__N_2493[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i9_3_lut_4_lut.init = 16'hf1e0;
    FD1P3IX spi_data__i21 (.D(wb_dat_o[5]), .SP(clk_enable_569), .CD(n6196), 
            .CK(clk), .Q(\spi_data[21] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i21.GSR = "ENABLED";
    FD1P3IX spi_data__i20 (.D(wb_dat_o[4]), .SP(clk_enable_569), .CD(n6196), 
            .CK(clk), .Q(\spi_data[20] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i20.GSR = "ENABLED";
    FD1P3IX spi_data__i19 (.D(wb_dat_o[3]), .SP(clk_enable_569), .CD(n6196), 
            .CK(clk), .Q(\spi_data[19] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i19.GSR = "ENABLED";
    FD1P3IX spi_data__i18 (.D(wb_dat_o[2]), .SP(clk_enable_569), .CD(n6196), 
            .CK(clk), .Q(\spi_data[18] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i18.GSR = "ENABLED";
    FD1P3IX spi_data__i17 (.D(wb_dat_o[1]), .SP(clk_enable_569), .CD(n6196), 
            .CK(clk), .Q(\spi_data[17] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i17.GSR = "ENABLED";
    LUT4 mux_428_i8_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[7]), 
         .D(quad_count_adj_324[7]), .Z(\spi_data_out_r_39__N_2493[7] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i8_3_lut_4_lut.init = 16'hf1e0;
    FD1P3IX spi_data__i16 (.D(wb_dat_o[0]), .SP(clk_enable_569), .CD(n6196), 
            .CK(clk), .Q(\spi_data[16] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i16.GSR = "ENABLED";
    FD1P3IX spi_data__i15 (.D(wb_dat_o[7]), .SP(clk_enable_577), .CD(n6196), 
            .CK(clk), .Q(\spi_data[15] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i15.GSR = "ENABLED";
    FD1P3IX spi_data__i14 (.D(wb_dat_o[6]), .SP(clk_enable_577), .CD(n6196), 
            .CK(clk), .Q(\spi_data[14] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i14.GSR = "ENABLED";
    FD1P3IX spi_data__i13 (.D(wb_dat_o[5]), .SP(clk_enable_577), .CD(n6196), 
            .CK(clk), .Q(\spi_data[13] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i13.GSR = "ENABLED";
    FD1P3IX spi_data__i12 (.D(wb_dat_o[4]), .SP(clk_enable_577), .CD(n6196), 
            .CK(clk), .Q(\spi_data[12] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i12.GSR = "ENABLED";
    FD1P3IX spi_data__i11 (.D(wb_dat_o[3]), .SP(clk_enable_577), .CD(n6196), 
            .CK(clk), .Q(\spi_data[11] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i11.GSR = "ENABLED";
    FD1P3IX spi_data__i10 (.D(wb_dat_o[2]), .SP(clk_enable_577), .CD(n6196), 
            .CK(clk), .Q(\spi_data[10] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i10.GSR = "ENABLED";
    FD1P3IX spi_data__i9 (.D(wb_dat_o[1]), .SP(clk_enable_577), .CD(n6196), 
            .CK(clk), .Q(\spi_data[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i9.GSR = "ENABLED";
    FD1P3IX spi_data__i8 (.D(wb_dat_o[0]), .SP(clk_enable_577), .CD(n6196), 
            .CK(clk), .Q(\spi_data[8] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i8.GSR = "ENABLED";
    FD1P3IX spi_data__i7 (.D(wb_dat_o[7]), .SP(clk_enable_584), .CD(n6196), 
            .CK(clk), .Q(\spi_data[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i7.GSR = "ENABLED";
    FD1P3IX spi_data__i6 (.D(wb_dat_o[6]), .SP(clk_enable_584), .CD(n6196), 
            .CK(clk), .Q(\spi_data[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i6.GSR = "ENABLED";
    FD1P3IX spi_data__i5 (.D(wb_dat_o[5]), .SP(clk_enable_584), .CD(n6196), 
            .CK(clk), .Q(\spi_data[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i5.GSR = "ENABLED";
    FD1P3IX spi_data__i4 (.D(wb_dat_o[4]), .SP(clk_enable_584), .CD(n6196), 
            .CK(clk), .Q(\spi_data[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i4.GSR = "ENABLED";
    FD1P3IX spi_data__i3 (.D(wb_dat_o[3]), .SP(clk_enable_584), .CD(n6196), 
            .CK(clk), .Q(\spi_data[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i3.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_757 (.A(spi_cmd[7]), .B(spi_cmd[15]), .Z(n30157)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_rep_757.init = 16'h4444;
    LUT4 mux_422_i10_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[9]), 
         .D(quad_count[9]), .Z(\spi_data_out_r_39__N_1083[9] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i10_3_lut_4_lut.init = 16'hf1e0;
    FD1P3IX spi_data__i2 (.D(wb_dat_o[2]), .SP(clk_enable_584), .CD(n6196), 
            .CK(clk), .Q(\spi_data[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i2.GSR = "ENABLED";
    FD1P3IX spi_data__i1 (.D(wb_dat_o[1]), .SP(clk_enable_584), .CD(n6196), 
            .CK(clk), .Q(\spi_data[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i1.GSR = "ENABLED";
    LUT4 mux_422_i9_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[8]), 
         .D(quad_count[8]), .Z(\spi_data_out_r_39__N_1083[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_4_lut_adj_606 (.A(spi_cmd[7]), .B(spi_cmd[15]), .C(n30158), 
         .D(n30194), .Z(n27197)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_3_lut_4_lut_adj_606.init = 16'h0004;
    LUT4 mux_428_i7_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[6]), 
         .D(quad_count_adj_324[6]), .Z(\spi_data_out_r_39__N_2493[6] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i6_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[5]), 
         .D(quad_count_adj_324[5]), .Z(\spi_data_out_r_39__N_2493[5] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i5_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[4]), 
         .D(quad_count_adj_324[4]), .Z(\spi_data_out_r_39__N_2493[4] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i4_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[3]), 
         .D(quad_count_adj_324[3]), .Z(\spi_data_out_r_39__N_2493[3] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i3_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[2]), 
         .D(quad_count_adj_324[2]), .Z(\spi_data_out_r_39__N_2493[2] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i2_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[1]), 
         .D(quad_count_adj_324[1]), .Z(\spi_data_out_r_39__N_2493[1] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_758 (.A(spi_addr[2]), .B(spi_cmd[2]), .Z(n30158)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_rep_758.init = 16'heeee;
    LUT4 mux_426_i21_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[20]), 
         .D(quad_count_adj_322[20]), .Z(\spi_data_out_r_39__N_2023[20] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i1_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[0]), 
         .D(quad_count_adj_326[0]), .Z(\spi_data_out_r_39__N_2258[0] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i32_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[31]), 
         .D(quad_count_adj_326[31]), .Z(\spi_data_out_r_39__N_2258[31] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i31_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[30]), 
         .D(quad_count_adj_326[30]), .Z(\spi_data_out_r_39__N_2258[30] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i30_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[29]), 
         .D(quad_count_adj_326[29]), .Z(\spi_data_out_r_39__N_2258[29] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i29_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[28]), 
         .D(quad_count_adj_326[28]), .Z(\spi_data_out_r_39__N_2258[28] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i28_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[27]), 
         .D(quad_count_adj_326[27]), .Z(\spi_data_out_r_39__N_2258[27] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i27_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[26]), 
         .D(quad_count_adj_326[26]), .Z(\spi_data_out_r_39__N_2258[26] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i14075_3_lut_3_lut_4_lut (.A(n30169), .B(spi_idle), .C(\address_7__N_549[1] ), 
         .D(wb_dat_o[3]), .Z(rd_en_N_717)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:73])
    defparam i14075_3_lut_3_lut_4_lut.init = 16'hf010;
    LUT4 i1_4_lut_adj_607 (.A(n1220[2]), .B(n26715), .C(spi_cmd_start_reg_N_745), 
         .D(n1220[4]), .Z(n26721)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_607.init = 16'h0004;
    LUT4 i1_4_lut_adj_608 (.A(n28290), .B(n30147), .C(n26771), .D(spi_addr[2]), 
         .Z(n26779)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_adj_608.init = 16'h0040;
    LUT4 mux_427_i26_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[25]), 
         .D(quad_count_adj_326[25]), .Z(\spi_data_out_r_39__N_2258[25] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i25_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[24]), 
         .D(quad_count_adj_326[24]), .Z(\spi_data_out_r_39__N_2258[24] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_422_i23_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[22]), 
         .D(quad_count[22]), .Z(\spi_data_out_r_39__N_1083[22] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_4_lut_adj_609 (.A(spi_addr[2]), .B(spi_cmd[2]), .C(spi_cmd[7]), 
         .D(n30194), .Z(n26641)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_3_lut_4_lut_adj_609.init = 16'hfffe;
    LUT4 mux_427_i24_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[23]), 
         .D(quad_count_adj_326[23]), .Z(\spi_data_out_r_39__N_2258[23] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i23_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[22]), 
         .D(quad_count_adj_326[22]), .Z(\spi_data_out_r_39__N_2258[22] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i22_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[21]), 
         .D(quad_count_adj_326[21]), .Z(\spi_data_out_r_39__N_2258[21] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i21_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[20]), 
         .D(quad_count_adj_326[20]), .Z(\spi_data_out_r_39__N_2258[20] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i20_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[19]), 
         .D(quad_count_adj_326[19]), .Z(\spi_data_out_r_39__N_2258[19] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17483_2_lut (.A(spi_byte_cnt[1]), .B(spi_byte_cnt[0]), .Z(n21[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/spi_ctrl.v(383[46:62])
    defparam i17483_2_lut.init = 16'h6666;
    LUT4 mux_427_i19_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[18]), 
         .D(quad_count_adj_326[18]), .Z(\spi_data_out_r_39__N_2258[18] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_610 (.A(n26655), .B(n30198), .C(n30154), .D(n27065), 
         .Z(n47_adj_203)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_610.init = 16'hffef;
    LUT4 mux_427_i18_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[17]), 
         .D(quad_count_adj_326[17]), .Z(\spi_data_out_r_39__N_2258[17] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_611 (.A(n30194), .B(n30084), .C(n30145), .D(n27057), 
         .Z(n27065)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_611.init = 16'hfffe;
    LUT4 i1_2_lut_adj_612 (.A(spi_addr[1]), .B(spi_addr[0]), .Z(n27057)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_adj_612.init = 16'heeee;
    LUT4 mux_427_i17_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[16]), 
         .D(quad_count_adj_326[16]), .Z(\spi_data_out_r_39__N_2258[16] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i16_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[15]), 
         .D(quad_count_adj_326[15]), .Z(\spi_data_out_r_39__N_2258[15] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i16_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX wr_data_i0_i1 (.D(n672[1]), .SP(clk_enable_756), .CK(clk), 
            .Q(wr_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i1.GSR = "ENABLED";
    LUT4 mux_427_i15_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[14]), 
         .D(quad_count_adj_326[14]), .Z(\spi_data_out_r_39__N_2258[14] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i14_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[13]), 
         .D(quad_count_adj_326[13]), .Z(\spi_data_out_r_39__N_2258[13] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i14_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX wr_data_i0_i2 (.D(n672[2]), .SP(clk_enable_756), .CK(clk), 
            .Q(wr_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i2.GSR = "ENABLED";
    FD1P3AX wr_data_i0_i3 (.D(n672[3]), .SP(clk_enable_756), .CK(clk), 
            .Q(wr_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i3.GSR = "ENABLED";
    FD1P3AX wr_data_i0_i4 (.D(n672[4]), .SP(clk_enable_756), .CK(clk), 
            .Q(wr_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i4.GSR = "ENABLED";
    FD1P3AX wr_data_i0_i5 (.D(n672[5]), .SP(clk_enable_756), .CK(clk), 
            .Q(wr_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i5.GSR = "ENABLED";
    FD1P3AX wr_data_i0_i6 (.D(n672[6]), .SP(clk_enable_756), .CK(clk), 
            .Q(wr_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i6.GSR = "ENABLED";
    FD1P3AX wr_data_i0_i7 (.D(n672[7]), .SP(clk_enable_756), .CK(clk), 
            .Q(wr_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i7.GSR = "ENABLED";
    LUT4 mux_427_i13_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[12]), 
         .D(quad_count_adj_326[12]), .Z(\spi_data_out_r_39__N_2258[12] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i12_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[11]), 
         .D(quad_count_adj_326[11]), .Z(\spi_data_out_r_39__N_2258[11] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i11_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[10]), 
         .D(quad_count_adj_326[10]), .Z(\spi_data_out_r_39__N_2258[10] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i10_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[9]), 
         .D(quad_count_adj_326[9]), .Z(\spi_data_out_r_39__N_2258[9] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_759 (.A(spi_addr[0]), .B(spi_addr[2]), .Z(n30159)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_759.init = 16'heeee;
    LUT4 i1_2_lut_rep_760 (.A(spi_addr[0]), .B(spi_cmd[0]), .Z(n30160)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_760.init = 16'heeee;
    LUT4 i1_2_lut_rep_669_3_lut (.A(spi_addr[0]), .B(spi_cmd[0]), .C(spi_addr[1]), 
         .Z(n30069)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_669_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_619_3_lut_4_lut (.A(spi_addr[0]), .B(spi_cmd[0]), 
         .C(spi_cmd[2]), .D(spi_addr[1]), .Z(n30019)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_619_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut_adj_613 (.A(spi_addr[0]), .B(spi_cmd[0]), .C(spi_addr[1]), 
         .D(n32), .Z(n27215)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_3_lut_4_lut_adj_613.init = 16'h0010;
    LUT4 mem_addr_1792_mux_6_i3_3_lut_4_lut (.A(n31067), .B(n30173), .C(n37[2]), 
         .D(wb_dat_o[2]), .Z(n2[2])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam mem_addr_1792_mux_6_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_614 (.A(n27037), .B(n26655), .C(n30154), .D(n27027), 
         .Z(n47_adj_204)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_614.init = 16'hffef;
    LUT4 mux_427_i9_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[8]), 
         .D(quad_count_adj_326[8]), .Z(\spi_data_out_r_39__N_2258[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_615 (.A(n26355), .B(n30198), .C(n30026), .D(n32), 
         .Z(n16815)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_615.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_616 (.A(spi_addr[0]), .B(spi_cmd[0]), .C(spi_cmd[7]), 
         .Z(n27077)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_3_lut_adj_616.init = 16'hfefe;
    LUT4 mem_addr_1792_mux_6_i6_3_lut_4_lut (.A(n31067), .B(n30173), .C(n37[5]), 
         .D(wb_dat_o[5]), .Z(n2[5])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam mem_addr_1792_mux_6_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut_adj_617 (.A(n30084), .B(n30157), .C(n30101), .D(spi_cmd[2]), 
         .Z(n27171)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_617.init = 16'h0004;
    LUT4 i1_2_lut_rep_756 (.A(spi_addr[0]), .B(spi_addr[1]), .Z(n30156)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_2_lut_rep_756.init = 16'h8888;
    LUT4 mem_addr_1792_mux_6_i2_3_lut_4_lut (.A(n31067), .B(n30173), .C(n37[1]), 
         .D(wb_dat_o[1]), .Z(n2[1])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam mem_addr_1792_mux_6_i2_3_lut_4_lut.init = 16'hf780;
    FD1S3AX address_i2 (.D(address_7__N_359[1]), .CK(clk), .Q(\address[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam address_i2.GSR = "ENABLED";
    FD1P3AY spi_cmd_i0_i1 (.D(wb_dat_o[1]), .SP(clk_enable_859), .CK(clk), 
            .Q(spi_cmd[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_761 (.A(spi_cmd[7]), .B(spi_addr[2]), .Z(n30161)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_rep_761.init = 16'heeee;
    LUT4 mux_427_i8_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[7]), 
         .D(quad_count_adj_326[7]), .Z(\spi_data_out_r_39__N_2258[7] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24160_4_lut (.A(spi_cmd_start_reg_N_745), .B(n1220[10]), .C(n1220[9]), 
         .D(n30136), .Z(n28573)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i24160_4_lut.init = 16'habaa;
    LUT4 i1_3_lut_rep_627_4_lut (.A(spi_cmd[7]), .B(spi_addr[2]), .C(n30084), 
         .D(n30194), .Z(n30027)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_3_lut_rep_627_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_618 (.A(mem_burst_cnt[3]), .B(mem_burst_cnt[7]), .C(mem_burst_cnt[6]), 
         .D(mem_burst_cnt[5]), .Z(n23343)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(355[47:82])
    defparam i1_4_lut_adj_618.init = 16'hfffe;
    LUT4 mem_addr_1792_mux_6_i8_3_lut_4_lut (.A(n31067), .B(n30173), .C(n37[7]), 
         .D(wb_dat_o[7]), .Z(n2[7])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam mem_addr_1792_mux_6_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 i13910_2_lut (.A(mem_burst_cnt[0]), .B(mem_burst_cnt[2]), .Z(n18233)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13910_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_619 (.A(n27089), .B(n30198), .C(n27081), .D(spi_cmd[15]), 
         .Z(n47_adj_205)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_619.init = 16'hfeff;
    LUT4 mux_427_i7_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[6]), 
         .D(quad_count_adj_326[6]), .Z(\spi_data_out_r_39__N_2258[6] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i6_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[5]), 
         .D(quad_count_adj_326[5]), .Z(\spi_data_out_r_39__N_2258[5] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i5_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[4]), 
         .D(quad_count_adj_326[4]), .Z(\spi_data_out_r_39__N_2258[4] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_620 (.A(n27177), .B(n32), .C(n30194), .D(n27077), 
         .Z(n27089)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_620.init = 16'hfffd;
    LUT4 mem_addr_1792_mux_6_i5_3_lut_4_lut (.A(n31067), .B(n30173), .C(n37[4]), 
         .D(wb_dat_o[4]), .Z(n2[4])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam mem_addr_1792_mux_6_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_adj_621 (.A(spi_addr[2]), .B(spi_cmd[2]), .Z(n27177)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_621.init = 16'h8888;
    LUT4 i398_2_lut_rep_818 (.A(n1220[9]), .B(mem_rdata_update_N_729), .Z(n31067)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i398_2_lut_rep_818.init = 16'heeee;
    LUT4 mem_addr_1792_mux_6_i4_3_lut_4_lut (.A(n31067), .B(n30173), .C(n37[3]), 
         .D(wb_dat_o[3]), .Z(n2[3])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam mem_addr_1792_mux_6_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_427_i4_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[3]), 
         .D(quad_count_adj_326[3]), .Z(\spi_data_out_r_39__N_2258[3] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_422_i18_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[17]), 
         .D(quad_count[17]), .Z(\spi_data_out_r_39__N_1083[17] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mem_addr_1792_mux_6_i1_3_lut_4_lut (.A(n31067), .B(n30173), .C(n37[0]), 
         .D(wb_dat_o[0]), .Z(n2[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam mem_addr_1792_mux_6_i1_3_lut_4_lut.init = 16'hf780;
    LUT4 mem_addr_1792_mux_6_i7_3_lut_4_lut (.A(n31067), .B(n30173), .C(n37[6]), 
         .D(wb_dat_o[6]), .Z(n2[6])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam mem_addr_1792_mux_6_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 mux_427_i3_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[2]), 
         .D(quad_count_adj_326[2]), .Z(\spi_data_out_r_39__N_2258[2] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_426_i20_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[19]), 
         .D(quad_count_adj_322[19]), .Z(\spi_data_out_r_39__N_2023[19] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_427_i2_3_lut_4_lut (.A(n26483), .B(n30096), .C(quad_buffer_adj_325[1]), 
         .D(quad_count_adj_326[1]), .Z(\spi_data_out_r_39__N_2258[1] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_427_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i1_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[4] ), 
         .D(\SLO_buf[14] ), .Z(\spi_data_out_r_39__N_5105[0] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i1_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i7413 (.BLUT(n23208), .ALUT(wr_en_N_701), .C0(n30136), .Z(n11758));
    LUT4 mux_158_i36_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[3] ), 
         .D(\SLO_buf[9] ), .Z(\spi_data_out_r_39__N_5105[35] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i36_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i24109_2_lut_3_lut_3_lut_4_lut (.A(n1220[9]), .B(mem_rdata_update_N_729), 
         .C(\address_7__N_549[1] ), .D(spi_addr_valid_N_732), .Z(n12446)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i24109_2_lut_3_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 mux_158_i35_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[2] ), 
         .D(\SLO_buf[8] ), .Z(\spi_data_out_r_39__N_5105[34] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i35_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i24178_4_lut_4_lut_rep_676 (.A(n31067), .B(n30173), .C(spi_addr_valid_N_732), 
         .D(\address_7__N_549[1] ), .Z(clk_enable_915)) /* synthesis lut_function=(A (B)+!A (C (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i24178_4_lut_4_lut_rep_676.init = 16'hd888;
    LUT4 mux_158_i34_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[1] ), 
         .D(\SLO_buf[7] ), .Z(\spi_data_out_r_39__N_5105[33] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i34_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_424_i1_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[0]), 
         .D(quad_count_adj_328[0]), .Z(\spi_data_out_r_39__N_1553[0] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i32_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[31]), 
         .D(quad_count_adj_328[31]), .Z(\spi_data_out_r_39__N_1553[31] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i33_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[0] ), 
         .D(\SLO_buf[6] ), .Z(\spi_data_out_r_39__N_5105[32] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i33_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_158_i16_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[19] ), 
         .D(\SLO_buf[29] ), .Z(\spi_data_out_r_39__N_5105[15] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i16_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_424_i31_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[30]), 
         .D(quad_count_adj_328[30]), .Z(\spi_data_out_r_39__N_1553[30] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i30_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[29]), 
         .D(quad_count_adj_328[29]), .Z(\spi_data_out_r_39__N_1553[29] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i29_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[28]), 
         .D(quad_count_adj_328[28]), .Z(\spi_data_out_r_39__N_1553[28] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i28_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[27]), 
         .D(quad_count_adj_328[27]), .Z(\spi_data_out_r_39__N_1553[27] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i15_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[18] ), 
         .D(\SLO_buf[28] ), .Z(\spi_data_out_r_39__N_5105[14] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i15_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_424_i27_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[26]), 
         .D(quad_count_adj_328[26]), .Z(\spi_data_out_r_39__N_1553[26] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i27_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX spi_cmd_i0_i2 (.D(wb_dat_o[2]), .SP(clk_enable_859), .CK(clk), 
            .Q(spi_cmd[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i2.GSR = "ENABLED";
    FD1P3AY spi_cmd_i0_i3 (.D(wb_dat_o[3]), .SP(clk_enable_859), .CK(clk), 
            .Q(spi_cmd[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i3.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i4 (.D(wb_dat_o[4]), .SP(clk_enable_859), .CK(clk), 
            .Q(spi_cmd[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i4.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i5 (.D(wb_dat_o[5]), .SP(clk_enable_859), .CK(clk), 
            .Q(spi_cmd[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i5.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i6 (.D(wb_dat_o[6]), .SP(clk_enable_859), .CK(clk), 
            .Q(spi_cmd[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i6.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i7 (.D(wb_dat_o[7]), .SP(clk_enable_859), .CK(clk), 
            .Q(spi_cmd[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i7.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i8 (.D(wb_dat_o[0]), .SP(clk_enable_867), .CK(clk), 
            .Q(spi_cmd[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i8.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i9 (.D(wb_dat_o[1]), .SP(clk_enable_867), .CK(clk), 
            .Q(spi_cmd[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i9.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i10 (.D(wb_dat_o[2]), .SP(clk_enable_867), .CK(clk), 
            .Q(spi_cmd[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i10.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i11 (.D(wb_dat_o[3]), .SP(clk_enable_867), .CK(clk), 
            .Q(spi_cmd[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i11.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i12 (.D(wb_dat_o[4]), .SP(clk_enable_867), .CK(clk), 
            .Q(spi_cmd[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i12.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i13 (.D(wb_dat_o[5]), .SP(clk_enable_867), .CK(clk), 
            .Q(spi_cmd[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i13.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i14 (.D(wb_dat_o[6]), .SP(clk_enable_867), .CK(clk), 
            .Q(spi_cmd[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i14.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i15 (.D(wb_dat_o[7]), .SP(clk_enable_867), .CK(clk), 
            .Q(spi_cmd[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i15.GSR = "ENABLED";
    LUT4 mux_158_i14_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[17] ), 
         .D(\SLO_buf[27] ), .Z(\spi_data_out_r_39__N_5105[13] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i14_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_426_i26_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[25]), 
         .D(quad_count_adj_322[25]), .Z(\spi_data_out_r_39__N_2023[25] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i26_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[25]), 
         .D(quad_count_adj_328[25]), .Z(\spi_data_out_r_39__N_1553[25] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i25_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[24]), 
         .D(quad_count_adj_328[24]), .Z(\spi_data_out_r_39__N_1553[24] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_adj_622 (.A(wr_en), .B(wb_sm), .Z(wb_we_i_N_344)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_adj_622.init = 16'h2222;
    LUT4 mux_158_i13_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[16] ), 
         .D(\SLO_buf[26] ), .Z(\spi_data_out_r_39__N_5105[12] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i13_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_424_i24_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[23]), 
         .D(quad_count_adj_328[23]), .Z(\spi_data_out_r_39__N_1553[23] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i12_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[15] ), 
         .D(\SLO_buf[25] ), .Z(\spi_data_out_r_39__N_5105[11] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i12_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_158_i11_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[14] ), 
         .D(\SLO_buf[24] ), .Z(\spi_data_out_r_39__N_5105[10] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i11_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i7814_3_lut (.A(spi_cmd_start_reg_N_745), .B(spi_idle_N_747), .C(spi_idle), 
         .Z(n12176)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(130[11] 133[31])
    defparam i7814_3_lut.init = 16'hdcdc;
    LUT4 mux_424_i23_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[22]), 
         .D(quad_count_adj_328[22]), .Z(\spi_data_out_r_39__N_1553[22] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i10_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[13] ), 
         .D(\SLO_buf[23] ), .Z(\spi_data_out_r_39__N_5105[9] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i10_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i7414_4_lut (.A(n28534), .B(spi_addr_valid_N_732), .C(n25421), 
         .D(n12), .Z(n11759)) /* synthesis lut_function=(A (B)+!A (B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i7414_4_lut.init = 16'hdddc;
    LUT4 i1_4_lut_adj_623 (.A(spi_idle), .B(n30169), .C(wb_dat_o[4]), 
         .D(wb_dat_o[3]), .Z(n23860)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:73])
    defparam i1_4_lut_adj_623.init = 16'hfffe;
    LUT4 mux_424_i22_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[21]), 
         .D(quad_count_adj_328[21]), .Z(\spi_data_out_r_39__N_1553[21] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23832_4_lut (.A(\address_7__N_549[1] ), .B(n28508), .C(n10254), 
         .D(n10255), .Z(n28534)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;
    defparam i23832_4_lut.init = 16'heeec;
    LUT4 mux_424_i21_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[20]), 
         .D(quad_count_adj_328[20]), .Z(\spi_data_out_r_39__N_1553[20] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23806_4_lut (.A(n1220[11]), .B(n28426), .C(n7970), .D(\address_7__N_549[1] ), 
         .Z(n28508)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i23806_4_lut.init = 16'heccc;
    LUT4 i1_4_lut_adj_624 (.A(n24183), .B(n1220[9]), .C(n6), .D(n30217), 
         .Z(n12)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_624.init = 16'ha0a8;
    LUT4 mux_424_i20_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[19]), 
         .D(quad_count_adj_328[19]), .Z(\spi_data_out_r_39__N_1553[19] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_1235_i1_3_lut (.A(n11758), .B(\address_7__N_549[1] ), .C(spi_cmd_start_reg_N_746), 
         .Z(wr_en_N_697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam mux_1235_i1_3_lut.init = 16'hcaca;
    LUT4 i1441_2_lut (.A(spi_cmd_cnt), .B(n1220[5]), .Z(spi_cmd_cnt_N_749)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1441_2_lut.init = 16'h6666;
    LUT4 mux_424_i19_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[18]), 
         .D(quad_count_adj_328[18]), .Z(\spi_data_out_r_39__N_1553[18] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i18_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[17]), 
         .D(quad_count_adj_328[17]), .Z(\spi_data_out_r_39__N_1553[17] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i17_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[16]), 
         .D(quad_count_adj_328[16]), .Z(\spi_data_out_r_39__N_1553[16] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_422_i17_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[16]), 
         .D(quad_count[16]), .Z(\spi_data_out_r_39__N_1083[16] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i16_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[15]), 
         .D(quad_count_adj_328[15]), .Z(\spi_data_out_r_39__N_1553[15] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i15_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[14]), 
         .D(quad_count_adj_328[14]), .Z(\spi_data_out_r_39__N_1553[14] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i14_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[13]), 
         .D(quad_count_adj_328[13]), .Z(\spi_data_out_r_39__N_1553[13] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_422_i16_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[15]), 
         .D(quad_count[15]), .Z(\spi_data_out_r_39__N_1083[15] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i16_3_lut_4_lut.init = 16'hf1e0;
    CCU2D mem_addr_1792_add_4_9 (.A0(spi_addr[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21900), .S0(n37[7]));   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_1792_add_4_9.INIT0 = 16'hfaaa;
    defparam mem_addr_1792_add_4_9.INIT1 = 16'h0000;
    defparam mem_addr_1792_add_4_9.INJECT1_0 = "NO";
    defparam mem_addr_1792_add_4_9.INJECT1_1 = "NO";
    CCU2D mem_addr_1792_add_4_7 (.A0(spi_addr[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_addr[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21899), .COUT(n21900), .S0(n37[5]), .S1(n37[6]));   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_1792_add_4_7.INIT0 = 16'hfaaa;
    defparam mem_addr_1792_add_4_7.INIT1 = 16'hfaaa;
    defparam mem_addr_1792_add_4_7.INJECT1_0 = "NO";
    defparam mem_addr_1792_add_4_7.INJECT1_1 = "NO";
    CCU2D mem_addr_1792_add_4_5 (.A0(spi_addr[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_addr[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21898), .COUT(n21899), .S0(n37[3]), .S1(n37[4]));   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_1792_add_4_5.INIT0 = 16'hfaaa;
    defparam mem_addr_1792_add_4_5.INIT1 = 16'hfaaa;
    defparam mem_addr_1792_add_4_5.INJECT1_0 = "NO";
    defparam mem_addr_1792_add_4_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(n30193), .B(spi_cmd[5]), .C(spi_cmd[9]), .D(n30093), 
         .Z(n26653)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_4_lut.init = 16'hfffe;
    CCU2D mem_addr_1792_add_4_3 (.A0(spi_addr[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_addr[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21897), .COUT(n21898), .S0(n37[1]), .S1(n37[2]));   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_1792_add_4_3.INIT0 = 16'hfaaa;
    defparam mem_addr_1792_add_4_3.INIT1 = 16'hfaaa;
    defparam mem_addr_1792_add_4_3.INJECT1_0 = "NO";
    defparam mem_addr_1792_add_4_3.INJECT1_1 = "NO";
    LUT4 mux_158_i9_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[12] ), 
         .D(\SLO_buf[22] ), .Z(\spi_data_out_r_39__N_5105[8] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i9_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_424_i13_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[12]), 
         .D(quad_count_adj_328[12]), .Z(\spi_data_out_r_39__N_1553[12] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_626_4_lut (.A(n30193), .B(spi_cmd[5]), .C(spi_cmd[9]), 
         .D(spi_cmd[0]), .Z(n30026)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_rep_626_4_lut.init = 16'hfeff;
    LUT4 i23588_2_lut_4_lut (.A(n30193), .B(spi_cmd[5]), .C(spi_cmd[9]), 
         .D(n30194), .Z(n28290)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i23588_2_lut_4_lut.init = 16'hfffe;
    LUT4 mux_158_i8_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[11] ), 
         .D(\SLO_buf[21] ), .Z(\spi_data_out_r_39__N_5105[7] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i8_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_424_i12_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[11]), 
         .D(quad_count_adj_328[11]), .Z(\spi_data_out_r_39__N_1553[11] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i7_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[10] ), 
         .D(\SLO_buf[20] ), .Z(\spi_data_out_r_39__N_5105[6] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i7_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_158_i6_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[9] ), 
         .D(\SLO_buf[19] ), .Z(\spi_data_out_r_39__N_5105[5] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i6_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_424_i11_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[10]), 
         .D(quad_count_adj_328[10]), .Z(\spi_data_out_r_39__N_1553[10] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_4_lut_adj_625 (.A(n30193), .B(spi_cmd[5]), .C(spi_cmd[9]), 
         .D(spi_addr[1]), .Z(n27081)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_4_lut_adj_625.init = 16'hfeff;
    CCU2D mem_addr_1792_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_addr[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n21897), .S1(n37[0]));   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_1792_add_4_1.INIT0 = 16'hF000;
    defparam mem_addr_1792_add_4_1.INIT1 = 16'h0555;
    defparam mem_addr_1792_add_4_1.INJECT1_0 = "NO";
    defparam mem_addr_1792_add_4_1.INJECT1_1 = "NO";
    LUT4 mux_158_i5_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[8] ), 
         .D(\SLO_buf[18] ), .Z(\spi_data_out_r_39__N_5105[4] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i5_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_424_i10_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[9]), 
         .D(quad_count_adj_328[9]), .Z(\spi_data_out_r_39__N_1553[9] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i9_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[8]), 
         .D(quad_count_adj_328[8]), .Z(\spi_data_out_r_39__N_1553[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i8_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[7]), 
         .D(quad_count_adj_328[7]), .Z(\spi_data_out_r_39__N_1553[7] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i7_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[6]), 
         .D(quad_count_adj_328[6]), .Z(\spi_data_out_r_39__N_1553[6] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i4_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[7] ), 
         .D(\SLO_buf[17] ), .Z(\spi_data_out_r_39__N_5105[3] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i4_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_424_i6_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[5]), 
         .D(quad_count_adj_328[5]), .Z(\spi_data_out_r_39__N_1553[5] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i5_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[4]), 
         .D(quad_count_adj_328[4]), .Z(\spi_data_out_r_39__N_1553[4] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i4_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[3]), 
         .D(quad_count_adj_328[3]), .Z(\spi_data_out_r_39__N_1553[3] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_426_i19_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[18]), 
         .D(quad_count_adj_322[18]), .Z(\spi_data_out_r_39__N_2023[18] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i3_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[2]), 
         .D(quad_count_adj_328[2]), .Z(\spi_data_out_r_39__N_1553[2] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_424_i2_3_lut_4_lut (.A(n16815), .B(n30159), .C(quad_buffer_adj_327[1]), 
         .D(quad_count_adj_328[1]), .Z(\spi_data_out_r_39__N_1553[1] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;
    defparam mux_424_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_4_lut_adj_626 (.A(n29997), .B(n30198), .C(spi_addr[2]), 
         .D(n30096), .Z(n47_adj_270)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_3_lut_4_lut_adj_626.init = 16'hfffe;
    LUT4 i1_2_lut_adj_627 (.A(spi_cmd_start_reg_N_745), .B(n1220[10]), .Z(n6196)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_adj_627.init = 16'h2222;
    LUT4 spi_cmd_start_I_15_2_lut_3_lut (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(spi_cmd_start_reg), .Z(spi_cmd_start)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(123[28:62])
    defparam spi_cmd_start_I_15_2_lut_3_lut.init = 16'hf2f2;
    LUT4 spi_xfer_done_I_10_2_lut_rep_769 (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .Z(n30169)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam spi_xfer_done_I_10_2_lut_rep_769.init = 16'h4444;
    LUT4 mux_158_i3_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[6] ), 
         .D(\SLO_buf[16] ), .Z(\spi_data_out_r_39__N_5105[2] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i3_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_158_i2_3_lut_4_lut (.A(n30156), .B(n16817), .C(\SLO_buf[5] ), 
         .D(\SLO_buf[15] ), .Z(\spi_data_out_r_39__N_5105[1] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mux_158_i2_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i1_2_lut_3_lut_4_lut_adj_628 (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(n1220[5]), .D(spi_idle), .Z(n23412)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B+((D)+!C)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam i1_2_lut_3_lut_4_lut_adj_628.init = 16'h00b0;
    LUT4 i24111_4_lut (.A(spi_byte_cnt[0]), .B(spi_byte_cnt[2]), .C(spi_byte_cnt[1]), 
         .D(spi_byte_cnt[3]), .Z(spi_data_valid_N_737)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/s_links/sources/spi_ctrl.v(331[12:16])
    defparam i24111_4_lut.init = 16'h0004;
    LUT4 i58_4_lut (.A(n29912), .B(spi_cmd_start), .C(spi_cmd_start_reg_N_745), 
         .D(n29), .Z(n32_adj_6711)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i58_4_lut.init = 16'hca0a;
    LUT4 i1_4_lut_adj_629 (.A(n24310), .B(n23469), .C(n26263), .D(n29997), 
         .Z(spi_data_out_r_39__N_2338)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_4_lut_adj_629.init = 16'h444c;
    LUT4 i1_3_lut (.A(spi_addr[0]), .B(n16815), .C(spi_addr[2]), .Z(n47_adj_271)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i1_3_lut.init = 16'hfdfd;
    LUT4 mux_422_i15_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[14]), 
         .D(quad_count[14]), .Z(\spi_data_out_r_39__N_1083[14] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_630 (.A(n26653), .B(n30198), .C(n26655), .D(spi_cmd[15]), 
         .Z(n24310)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_630.init = 16'hfeff;
    LUT4 i1_3_lut_rep_659_4_lut (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(wb_dat_o[3]), .D(spi_idle), .Z(n30059)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam i1_3_lut_rep_659_4_lut.init = 16'hfff4;
    LUT4 mux_422_i14_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[13]), 
         .D(quad_count[13]), .Z(\spi_data_out_r_39__N_1083[13] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i1_3_lut_4_lut_adj_631 (.A(n16817), .B(n30102), .C(\SLO_buf[4]_adj_272 ), 
         .D(\SLO_buf[14]_adj_273 ), .Z(\spi_data_out_r_39__N_4419[0] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i1_3_lut_4_lut_adj_631.init = 16'hf1e0;
    LUT4 i13054_2_lut_4_lut (.A(n23343), .B(n18233), .C(n30211), .D(mem_rdata[0]), 
         .Z(n672[0])) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(355[47:82])
    defparam i13054_2_lut_4_lut.init = 16'hff04;
    LUT4 i12910_2_lut_4_lut (.A(n23343), .B(n18233), .C(n30211), .D(mem_rdata[1]), 
         .Z(n672[1])) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(355[47:82])
    defparam i12910_2_lut_4_lut.init = 16'hff04;
    LUT4 i12901_2_lut_4_lut (.A(n23343), .B(n18233), .C(n30211), .D(mem_rdata[2]), 
         .Z(n672[2])) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(355[47:82])
    defparam i12901_2_lut_4_lut.init = 16'hff04;
    LUT4 mux_158_i36_3_lut_4_lut_adj_632 (.A(n16817), .B(n30102), .C(\SLO_buf[3]_adj_274 ), 
         .D(\SLO_buf[9]_adj_275 ), .Z(\spi_data_out_r_39__N_4419[35] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i36_3_lut_4_lut_adj_632.init = 16'hf1e0;
    LUT4 i12892_2_lut_4_lut (.A(n23343), .B(n18233), .C(n30211), .D(mem_rdata[3]), 
         .Z(n672[3])) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(355[47:82])
    defparam i12892_2_lut_4_lut.init = 16'hff04;
    LUT4 i1_4_lut_adj_633 (.A(n28290), .B(n30198), .C(n32), .D(n27127), 
         .Z(spi_data_out_r_39__N_4505)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_633.init = 16'h0100;
    LUT4 i1_4_lut_adj_634 (.A(n30197), .B(spi_cmd[7]), .C(spi_addr[2]), 
         .D(n30154), .Z(n27127)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_634.init = 16'h0200;
    LUT4 i1_3_lut_4_lut_adj_635 (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(wb_dat_o[4]), .D(spi_idle), .Z(n7970)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam i1_3_lut_4_lut_adj_635.init = 16'hfff4;
    LUT4 i12891_2_lut_4_lut (.A(n23343), .B(n18233), .C(n30211), .D(mem_rdata[4]), 
         .Z(n672[4])) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(355[47:82])
    defparam i12891_2_lut_4_lut.init = 16'hff04;
    LUT4 mux_426_i18_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[17]), 
         .D(quad_count_adj_322[17]), .Z(\spi_data_out_r_39__N_2023[17] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_426_i17_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[16]), 
         .D(quad_count_adj_322[16]), .Z(\spi_data_out_r_39__N_2023[16] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_4_lut_adj_636 (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(n30216), .D(spi_idle), .Z(n24198)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam i1_3_lut_4_lut_adj_636.init = 16'hfff4;
    LUT4 mux_422_i8_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[7]), 
         .D(quad_count[7]), .Z(\spi_data_out_r_39__N_1083[7] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_422_i7_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[6]), 
         .D(quad_count[6]), .Z(\spi_data_out_r_39__N_1083[6] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12888_2_lut_4_lut (.A(n23343), .B(n18233), .C(n30211), .D(mem_rdata[5]), 
         .Z(n672[5])) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(355[47:82])
    defparam i12888_2_lut_4_lut.init = 16'hff04;
    LUT4 mux_422_i21_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[20]), 
         .D(quad_count[20]), .Z(\spi_data_out_r_39__N_1083[20] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_426_i16_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[15]), 
         .D(quad_count_adj_322[15]), .Z(\spi_data_out_r_39__N_2023[15] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12879_2_lut_4_lut (.A(n23343), .B(n18233), .C(n30211), .D(mem_rdata[6]), 
         .Z(n672[6])) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(355[47:82])
    defparam i12879_2_lut_4_lut.init = 16'hff04;
    LUT4 i1_3_lut_adj_637 (.A(\status_cntr[12] ), .B(n29985), .C(resetn_c), 
         .Z(n25212)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_adj_637.init = 16'h4040;
    LUT4 mux_158_i35_3_lut_4_lut_adj_638 (.A(n16817), .B(n30102), .C(\SLO_buf[2]_adj_276 ), 
         .D(\SLO_buf[8]_adj_277 ), .Z(\spi_data_out_r_39__N_4419[34] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i35_3_lut_4_lut_adj_638.init = 16'hf1e0;
    LUT4 i24001_2_lut_3_lut_4_lut (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(\address_7__N_549[1] ), .D(spi_idle), .Z(n24183)) /* synthesis lut_function=(!(A (C (D))+!A (B (C)+!B (C (D))))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam i24001_2_lut_3_lut_4_lut.init = 16'h0fbf;
    LUT4 i1_2_lut_adj_639 (.A(spi_byte_cnt[1]), .B(n23360), .Z(clk_enable_561)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_639.init = 16'h4444;
    LUT4 mux_426_i15_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[14]), 
         .D(quad_count_adj_322[14]), .Z(\spi_data_out_r_39__N_2023[14] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i34_3_lut_4_lut_adj_640 (.A(n16817), .B(n30102), .C(\SLO_buf[1]_adj_278 ), 
         .D(\SLO_buf[7]_adj_279 ), .Z(\spi_data_out_r_39__N_4419[33] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i34_3_lut_4_lut_adj_640.init = 16'hf1e0;
    LUT4 mux_158_i33_3_lut_4_lut_adj_641 (.A(n16817), .B(n30102), .C(\SLO_buf[0]_adj_280 ), 
         .D(\SLO_buf[6]_adj_281 ), .Z(\spi_data_out_r_39__N_4419[32] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i33_3_lut_4_lut_adj_641.init = 16'hf1e0;
    LUT4 i12866_2_lut_4_lut (.A(n23343), .B(n18233), .C(n30211), .D(mem_rdata[7]), 
         .Z(n672[7])) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(355[47:82])
    defparam i12866_2_lut_4_lut.init = 16'hff04;
    LUT4 i1_4_lut_adj_642 (.A(spi_byte_cnt[3]), .B(n30054), .C(spi_byte_cnt[2]), 
         .D(spi_byte_cnt[0]), .Z(n23360)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_642.init = 16'h0400;
    LUT4 spi_xfer_done_I_0_240_2_lut_rep_674_3_lut (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(spi_idle), .Z(n30074)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam spi_xfer_done_I_0_240_2_lut_rep_674_3_lut.init = 16'hf4f4;
    LUT4 i1_4_lut_adj_643 (.A(n27215), .B(n30198), .C(n27211), .D(n30084), 
         .Z(clear_intrpt_N_3072)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_4_lut_adj_643.init = 16'h0020;
    LUT4 i1_4_lut_adj_644 (.A(n30194), .B(spi_cmd[7]), .C(spi_cmd[2]), 
         .D(n30195), .Z(n27211)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_644.init = 16'h0100;
    CCU2D mem_burst_cnt_1790_add_4_9 (.A0(mem_burst_cnt[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21890), .S0(n37_adj_7039[7]));   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_1790_add_4_9.INIT0 = 16'hfaaa;
    defparam mem_burst_cnt_1790_add_4_9.INIT1 = 16'h0000;
    defparam mem_burst_cnt_1790_add_4_9.INJECT1_0 = "NO";
    defparam mem_burst_cnt_1790_add_4_9.INJECT1_1 = "NO";
    LUT4 mux_426_i14_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[13]), 
         .D(quad_count_adj_322[13]), .Z(\spi_data_out_r_39__N_2023[13] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_adj_645 (.A(spi_byte_cnt[1]), .B(n23360), .Z(clk_enable_577)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_adj_645.init = 16'h8888;
    LUT4 mux_158_i16_3_lut_4_lut_adj_646 (.A(n16817), .B(n30102), .C(\SLO_buf[19]_adj_282 ), 
         .D(\SLO_buf[29]_adj_283 ), .Z(\spi_data_out_r_39__N_4419[15] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i16_3_lut_4_lut_adj_646.init = 16'hf1e0;
    LUT4 mux_422_i6_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[5]), 
         .D(quad_count[5]), .Z(\spi_data_out_r_39__N_1083[5] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i6_3_lut_4_lut.init = 16'hf1e0;
    CCU2D mem_burst_cnt_1790_add_4_7 (.A0(mem_burst_cnt[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(mem_burst_cnt[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n21889), .COUT(n21890), .S0(n37_adj_7039[5]), 
          .S1(n37_adj_7039[6]));   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_1790_add_4_7.INIT0 = 16'hfaaa;
    defparam mem_burst_cnt_1790_add_4_7.INIT1 = 16'hfaaa;
    defparam mem_burst_cnt_1790_add_4_7.INJECT1_0 = "NO";
    defparam mem_burst_cnt_1790_add_4_7.INJECT1_1 = "NO";
    CCU2D mem_burst_cnt_1790_add_4_5 (.A0(mem_burst_cnt[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(mem_burst_cnt[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n21888), .COUT(n21889), .S0(n37_adj_7039[3]), 
          .S1(n37_adj_7039[4]));   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_1790_add_4_5.INIT0 = 16'hfaaa;
    defparam mem_burst_cnt_1790_add_4_5.INIT1 = 16'hfaaa;
    defparam mem_burst_cnt_1790_add_4_5.INJECT1_0 = "NO";
    defparam mem_burst_cnt_1790_add_4_5.INJECT1_1 = "NO";
    CCU2D mem_burst_cnt_1790_add_4_3 (.A0(mem_burst_cnt[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(mem_burst_cnt[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n21887), .COUT(n21888), .S0(n37_adj_7039[1]), 
          .S1(n37_adj_7039[2]));   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_1790_add_4_3.INIT0 = 16'hfaaa;
    defparam mem_burst_cnt_1790_add_4_3.INIT1 = 16'hfaaa;
    defparam mem_burst_cnt_1790_add_4_3.INJECT1_0 = "NO";
    defparam mem_burst_cnt_1790_add_4_3.INJECT1_1 = "NO";
    CCU2D mem_burst_cnt_1790_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(mem_burst_cnt[0]), .B1(n18233), .C1(n30211), 
          .D1(n23343), .COUT(n21887), .S1(n37_adj_7039[0]));   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_1790_add_4_1.INIT0 = 16'hF000;
    defparam mem_burst_cnt_1790_add_4_1.INIT1 = 16'h5559;
    defparam mem_burst_cnt_1790_add_4_1.INJECT1_0 = "NO";
    defparam mem_burst_cnt_1790_add_4_1.INJECT1_1 = "NO";
    LUT4 mux_422_i5_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[4]), 
         .D(quad_count[4]), .Z(\spi_data_out_r_39__N_1083[4] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1478_3_lut_rep_773 (.A(mem_wr), .B(wr_en), .C(mem_rdata_update_N_729), 
         .Z(n30173)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1478_3_lut_rep_773.init = 16'hcaca;
    LUT4 i24114_2_lut_4_lut_4_lut_2_lut_3_lut (.A(n1220[9]), .B(mem_rdata_update_N_729), 
         .C(n1220[5]), .Z(n12460)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i24114_2_lut_4_lut_4_lut_2_lut_3_lut.init = 16'h1010;
    LUT4 mux_426_i13_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[12]), 
         .D(quad_count_adj_322[12]), .Z(\spi_data_out_r_39__N_2023[12] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_4_lut_adj_647 (.A(n30194), .B(n30196), .C(spi_addr[1]), 
         .D(spi_cmd[15]), .Z(n26355)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_3_lut_4_lut_adj_647.init = 16'hefff;
    LUT4 mux_158_i15_3_lut_4_lut_adj_648 (.A(n16817), .B(n30102), .C(\SLO_buf[18]_adj_284 ), 
         .D(\SLO_buf[28]_adj_285 ), .Z(\spi_data_out_r_39__N_4419[14] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i15_3_lut_4_lut_adj_648.init = 16'hf1e0;
    LUT4 i23742_3_lut_4_lut (.A(n1220[9]), .B(mem_rdata_update_N_729), .C(spi_addr_valid_N_732), 
         .D(n1220[6]), .Z(n28444)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i23742_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_158_i14_3_lut_4_lut_adj_649 (.A(n16817), .B(n30102), .C(\SLO_buf[17]_adj_286 ), 
         .D(\SLO_buf[27]_adj_287 ), .Z(\spi_data_out_r_39__N_4419[13] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i14_3_lut_4_lut_adj_649.init = 16'hf1e0;
    LUT4 mux_422_i13_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[12]), 
         .D(quad_count[12]), .Z(\spi_data_out_r_39__N_1083[12] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_650 (.A(n27229), .B(n30198), .C(n32), .D(n30084), 
         .Z(spi_data_out_r_39__N_4848)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_650.init = 16'h0002;
    LUT4 mux_422_i4_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[3]), 
         .D(quad_count[3]), .Z(\spi_data_out_r_39__N_1083[3] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_422_i3_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[2]), 
         .D(quad_count[2]), .Z(\spi_data_out_r_39__N_1083[2] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_651 (.A(n30194), .B(n27223), .C(spi_addr[2]), .D(spi_cmd[7]), 
         .Z(n27229)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_651.init = 16'h0004;
    LUT4 mux_426_i12_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[11]), 
         .D(quad_count_adj_322[11]), .Z(\spi_data_out_r_39__N_2023[11] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i13_3_lut_4_lut_adj_652 (.A(n16817), .B(n30102), .C(\SLO_buf[16]_adj_288 ), 
         .D(\SLO_buf[26]_adj_289 ), .Z(\spi_data_out_r_39__N_4419[12] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i13_3_lut_4_lut_adj_652.init = 16'hf1e0;
    LUT4 mux_426_i11_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[10]), 
         .D(quad_count_adj_322[10]), .Z(\spi_data_out_r_39__N_2023[10] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i24184_3_lut_rep_625_3_lut_4_lut (.A(n1220[9]), .B(mem_rdata_update_N_729), 
         .C(n1220[5]), .D(n30173), .Z(clk_enable_1128)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i24184_3_lut_rep_625_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_158_i12_3_lut_4_lut_adj_653 (.A(n16817), .B(n30102), .C(\SLO_buf[15]_adj_290 ), 
         .D(\SLO_buf[25]_adj_291 ), .Z(\spi_data_out_r_39__N_4419[11] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i12_3_lut_4_lut_adj_653.init = 16'hf1e0;
    LUT4 mux_158_i11_3_lut_4_lut_adj_654 (.A(n16817), .B(n30102), .C(\SLO_buf[14]_adj_273 ), 
         .D(\SLO_buf[24]_adj_292 ), .Z(\spi_data_out_r_39__N_4419[10] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i11_3_lut_4_lut_adj_654.init = 16'hf1e0;
    LUT4 mux_158_i10_3_lut_4_lut_adj_655 (.A(n16817), .B(n30102), .C(\SLO_buf[13]_adj_293 ), 
         .D(\SLO_buf[23]_adj_294 ), .Z(\spi_data_out_r_39__N_4419[9] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i10_3_lut_4_lut_adj_655.init = 16'hf1e0;
    LUT4 i2_1_lut_rep_782 (.A(spi_byte_cnt[0]), .Z(n30182)) /* synthesis lut_function=(!(A)) */ ;
    defparam i2_1_lut_rep_782.init = 16'h5555;
    LUT4 i1_3_lut_3_lut (.A(spi_byte_cnt[0]), .B(spi_byte_cnt[1]), .C(spi_byte_cnt[2]), 
         .Z(n27365)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_3_lut_3_lut.init = 16'h0404;
    LUT4 mux_158_i9_3_lut_4_lut_adj_656 (.A(n16817), .B(n30102), .C(\SLO_buf[12]_adj_295 ), 
         .D(\SLO_buf[22]_adj_296 ), .Z(\spi_data_out_r_39__N_4419[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i9_3_lut_4_lut_adj_656.init = 16'hf1e0;
    LUT4 resetn_I_0_1_lut_rep_785 (.A(resetn_c), .Z(n30185)) /* synthesis lut_function=(!(A)) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_I_0_1_lut_rep_785.init = 16'h5555;
    LUT4 reduce_or_1173_i1_4_lut_4_lut (.A(resetn_c), .B(n25885), .C(n30087), 
         .D(\quad_homing[1] ), .Z(n1)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam reduce_or_1173_i1_4_lut_4_lut.init = 16'h55d5;
    LUT4 i1_3_lut_3_lut_adj_657 (.A(resetn_c), .B(spi_sdo_valid), .C(mem_rdata_update), 
         .Z(clk_enable_963)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_3_lut_adj_657.init = 16'hfdfd;
    LUT4 i1_2_lut_rep_588_3_lut_3_lut (.A(resetn_c), .B(n30010), .C(\spi_addr_r[0] ), 
         .Z(clk_enable_686)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_rep_588_3_lut_3_lut.init = 16'h5d5d;
    LUT4 i1842_2_lut_4_lut_4_lut (.A(resetn_c), .B(spi_cmd_valid), .C(spi_scsn_dly), 
         .D(spi_scsn_c), .Z(clk_enable_776)) /* synthesis lut_function=((B+!(C+!(D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1842_2_lut_4_lut_4_lut.init = 16'hdfdd;
    LUT4 i2014_4_lut_4_lut (.A(resetn_c), .B(n26077), .C(n24066), .D(n30062), 
         .Z(clk_enable_260)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2014_4_lut_4_lut.init = 16'hd555;
    LUT4 resetn_N_2639_I_0_2_lut_2_lut (.A(resetn_c), .B(clear_intrpt), 
         .Z(intrpt_out_N_2642)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_N_2639_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 resetn_N_3065_I_0_2_lut_2_lut (.A(resetn_c), .B(clear_intrpt_adj_297), 
         .Z(intrpt_out_N_3068)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_N_3065_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1870_4_lut_4_lut (.A(resetn_c), .B(n28540), .C(n30035), .D(n23537), 
         .Z(clk_enable_263)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1870_4_lut_4_lut.init = 16'h7555;
    LUT4 i1854_2_lut_2_lut (.A(resetn_c), .B(quad_set_valid_N_1158), .Z(clk_enable_807)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1854_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_2_lut (.A(resetn_c), .B(n20598), .Z(n8400)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_2_lut.init = 16'hdddd;
    LUT4 i24155_4_lut_4_lut_4_lut (.A(resetn_c), .B(n12467), .C(n20647), 
         .D(n18654), .Z(n12435)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i24155_4_lut_4_lut_4_lut.init = 16'haa20;
    LUT4 i1_4_lut_4_lut_adj_658 (.A(resetn_c), .B(n4), .C(n30070), .D(n26873), 
         .Z(clk_enable_320)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_4_lut_adj_658.init = 16'h5d55;
    LUT4 reduce_or_1201_i1_4_lut_4_lut (.A(resetn_c), .B(n25877), .C(n30075), 
         .D(\quad_homing[1]_adj_298 ), .Z(n1_adj_299)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam reduce_or_1201_i1_4_lut_4_lut.init = 16'h55d5;
    LUT4 i1861_4_lut_4_lut (.A(resetn_c), .B(n30199), .C(n23916), .D(n26821), 
         .Z(clk_enable_684)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1861_4_lut_4_lut.init = 16'hd555;
    LUT4 i1_4_lut_4_lut_adj_659 (.A(resetn_c), .B(n26089), .C(n24066), 
         .D(n26091), .Z(clk_enable_255)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_4_lut_adj_659.init = 16'hd555;
    LUT4 i1_3_lut_4_lut_4_lut (.A(resetn_c), .B(EM_STOP), .C(clk_enable_259), 
         .D(n29996), .Z(clk_enable_23)) /* synthesis lut_function=((B ((D)+!C)+!B (D))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hff5d;
    LUT4 i2006_3_lut_3_lut (.A(resetn_c), .B(n23916), .C(n26947), .Z(clk_enable_253)) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2006_3_lut_3_lut.init = 16'hd5d5;
    LUT4 i1_3_lut_3_lut_adj_660 (.A(resetn_c), .B(pwm_out_N_3169), .C(pwm_out_N_3153), 
         .Z(clk_enable_15)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_3_lut_adj_660.init = 16'hfdfd;
    LUT4 i1_4_lut_4_lut_adj_661 (.A(resetn_c), .B(\spi_addr_r[7] ), .C(n26107), 
         .D(n30214), .Z(n26113)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_4_lut_adj_661.init = 16'hfffd;
    LUT4 resetn_N_2994_I_0_2_lut_2_lut (.A(resetn_c), .B(clear_intrpt_adj_300), 
         .Z(intrpt_out_N_2997)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_N_2994_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1859_4_lut_4_lut (.A(resetn_c), .B(n25993), .C(n24066), .D(n30062), 
         .Z(clk_enable_687)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1859_4_lut_4_lut.init = 16'hd555;
    LUT4 i1_2_lut_rep_589_4_lut_4_lut (.A(resetn_c), .B(n30045), .C(n28524), 
         .D(n23916), .Z(clk_enable_759)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_rep_589_4_lut_4_lut.init = 16'h5d55;
    LUT4 i1843_2_lut_4_lut_4_lut (.A(resetn_c), .B(clk_enable_48), .C(spi_scsn_dly), 
         .D(spi_scsn_c), .Z(clk_enable_624)) /* synthesis lut_function=(!(A (B (C+!(D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1843_2_lut_4_lut_4_lut.init = 16'h7f77;
    LUT4 i1860_2_lut_3_lut_4_lut_4_lut (.A(resetn_c), .B(n30033), .C(n23526), 
         .D(n30035), .Z(clk_enable_727)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1860_2_lut_3_lut_4_lut_4_lut.init = 16'hd555;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(resetn_c), .B(n11008), .C(pwm_out_1_N_6491), 
         .D(EM_STOP), .Z(clk_enable_613)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut_2_lut_adj_662 (.A(resetn_c), .B(spi_sdo_valid_N_296), 
         .Z(clk_enable_961)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_2_lut_adj_662.init = 16'hdddd;
    LUT4 i1855_4_lut_4_lut (.A(resetn_c), .B(n30011), .C(n26957), .D(n23916), 
         .Z(clk_enable_520)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1855_4_lut_4_lut.init = 16'hd555;
    LUT4 i1973_4_lut_4_lut (.A(resetn_c), .B(n28364), .C(n24065), .D(n26033), 
         .Z(clk_enable_232)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1973_4_lut_4_lut.init = 16'h7555;
    LUT4 i1_3_lut_4_lut_4_lut_adj_663 (.A(resetn_c), .B(EM_STOP), .C(clk_enable_254), 
         .D(n29995), .Z(clk_enable_28)) /* synthesis lut_function=((B ((D)+!C)+!B (D))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_663.init = 16'hff5d;
    LUT4 i1_4_lut_4_lut_adj_664 (.A(resetn_c), .B(n28514), .C(n23916), 
         .D(n26563), .Z(clk_enable_226)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_4_lut_adj_664.init = 16'h7555;
    LUT4 i1865_4_lut_4_lut (.A(resetn_c), .B(n30062), .C(n23916), .D(n26821), 
         .Z(clk_enable_639)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1865_4_lut_4_lut.init = 16'hd555;
    LUT4 i1845_2_lut_4_lut_4_lut (.A(resetn_c), .B(spi_cmd_valid), .C(spi_scsn_dly), 
         .D(spi_scsn_c), .Z(clk_enable_228)) /* synthesis lut_function=(!(A (B (C+!(D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1845_2_lut_4_lut_4_lut.init = 16'h7f77;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_665 (.A(resetn_c), .B(n11008), .C(pwm_out_3_N_6530), 
         .D(EM_STOP), .Z(clk_enable_1105)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_665.init = 16'hfff7;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_666 (.A(resetn_c), .B(n11008), .C(pwm_out_4_N_6549), 
         .D(EM_STOP), .Z(clk_enable_1107)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_666.init = 16'hfff7;
    LUT4 i1853_4_lut_4_lut (.A(resetn_c), .B(n26841), .C(n23916), .D(n26843), 
         .Z(clk_enable_757)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1853_4_lut_4_lut.init = 16'hd555;
    LUT4 i2002_4_lut_4_lut (.A(resetn_c), .B(n26023), .C(n24065), .D(n28366), 
         .Z(clk_enable_245)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2002_4_lut_4_lut.init = 16'h55d5;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_667 (.A(resetn_c), .B(n11008), .C(pwm_out_2_N_6511), 
         .D(EM_STOP), .Z(clk_enable_22)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_667.init = 16'hfff7;
    LUT4 i1_4_lut_4_lut_adj_668 (.A(resetn_c), .B(n23916), .C(n30022), 
         .D(n26415), .Z(clk_enable_488)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_4_lut_adj_668.init = 16'h5d55;
    LUT4 i1934_2_lut_4_lut_4_lut (.A(resetn_c), .B(n30199), .C(n23916), 
         .D(n26633), .Z(clk_enable_641)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1934_2_lut_4_lut_4_lut.init = 16'hd555;
    LUT4 i1869_4_lut_4_lut (.A(resetn_c), .B(n23537), .C(n30035), .D(n25833), 
         .Z(clk_enable_638)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1869_4_lut_4_lut.init = 16'hd555;
    LUT4 i1_2_lut_4_lut_4_lut (.A(resetn_c), .B(n30036), .C(n23916), .D(n26435), 
         .Z(clk_enable_959)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_4_lut_4_lut.init = 16'hd555;
    LUT4 i1_4_lut_4_lut_adj_669 (.A(resetn_c), .B(n18440), .C(n30035), 
         .D(n26249), .Z(clk_enable_235)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_4_lut_adj_669.init = 16'h7555;
    LUT4 resetn_N_2710_I_0_2_lut_2_lut (.A(resetn_c), .B(clear_intrpt_adj_301), 
         .Z(intrpt_out_N_2713)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_N_2710_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i75_2_lut_3_lut_3_lut (.A(resetn_c), .B(n11008), .C(EM_STOP), 
         .Z(n57)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i75_2_lut_3_lut_3_lut.init = 16'hfdfd;
    LUT4 i1878_2_lut_2_lut (.A(resetn_c), .B(reset_r_N_4129), .Z(clk_enable_761)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1878_2_lut_2_lut.init = 16'hdddd;
    LUT4 wb_rst_i_I_0_3_lut_rep_680_3_lut (.A(resetn_c), .B(spi_scsn_dly), 
         .C(spi_scsn_c), .Z(n30080)) /* synthesis lut_function=(!(A (B+!(C)))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam wb_rst_i_I_0_3_lut_rep_680_3_lut.init = 16'h7575;
    LUT4 i1_2_lut_rep_598_3_lut_3_lut (.A(resetn_c), .B(n11008), .C(EM_STOP), 
         .Z(n29998)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_rep_598_3_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_4_lut_4_lut_adj_670 (.A(resetn_c), .B(n28514), .C(n23916), 
         .D(n26539), .Z(clk_enable_738)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_4_lut_adj_670.init = 16'h7555;
    LUT4 reduce_or_1194_i1_4_lut_4_lut (.A(resetn_c), .B(n25881), .C(n30095), 
         .D(\quad_homing[1]_adj_302 ), .Z(n1_adj_303)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam reduce_or_1194_i1_4_lut_4_lut.init = 16'h55d5;
    LUT4 i1_4_lut_4_lut_adj_671 (.A(resetn_c), .B(n28516), .C(n23916), 
         .D(n26515), .Z(clk_enable_652)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_4_lut_adj_671.init = 16'h7555;
    LUT4 i1862_2_lut_2_lut (.A(resetn_c), .B(quad_set_valid_N_2098), .Z(clk_enable_683)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1862_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_672 (.A(resetn_c), .B(n30022), .C(n23526), 
         .D(n30035), .Z(clk_enable_211)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_672.init = 16'h7555;
    LUT4 i684_2_lut_2_lut (.A(resetn_c), .B(pwm_out_N_3169), .Z(n2109)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i684_2_lut_2_lut.init = 16'hdddd;
    LUT4 reduce_or_1180_i1_4_lut_4_lut (.A(resetn_c), .B(n25893), .C(n30055), 
         .D(\quad_homing[1]_adj_304 ), .Z(n1_adj_305)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam reduce_or_1180_i1_4_lut_4_lut.init = 16'h55d5;
    LUT4 reduce_or_1208_i1_4_lut_4_lut (.A(resetn_c), .B(n25869), .C(n30043), 
         .D(\quad_homing[1]_adj_306 ), .Z(n1_adj_307)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam reduce_or_1208_i1_4_lut_4_lut.init = 16'h55d5;
    LUT4 reduce_or_1187_i1_4_lut_4_lut (.A(resetn_c), .B(n25873), .C(n30091), 
         .D(\quad_homing[1]_adj_308 ), .Z(n1_adj_309)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam reduce_or_1187_i1_4_lut_4_lut.init = 16'h55d5;
    LUT4 i2018_4_lut_4_lut (.A(resetn_c), .B(n28476), .C(n24066), .D(n26059), 
         .Z(clk_enable_32)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2018_4_lut_4_lut.init = 16'h7555;
    LUT4 resetn_N_2852_I_0_2_lut_2_lut (.A(resetn_c), .B(clear_intrpt_adj_310), 
         .Z(intrpt_out_N_2855)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_N_2852_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_rep_587_3_lut_3_lut (.A(resetn_c), .B(n30010), .C(\spi_addr_r[0] ), 
         .Z(clk_enable_178)) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_rep_587_3_lut_3_lut.init = 16'hd5d5;
    LUT4 resetn_N_2781_I_0_2_lut_2_lut (.A(resetn_c), .B(clear_intrpt_adj_311), 
         .Z(intrpt_out_N_2784)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_N_2781_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1856_2_lut_2_lut (.A(resetn_c), .B(quad_set_valid_N_1393), .Z(clk_enable_842)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1856_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_673 (.A(resetn_c), .B(n18440), .C(n23916), 
         .D(n27013), .Z(clk_enable_627)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_673.init = 16'h7555;
    LUT4 i1970_4_lut_4_lut (.A(resetn_c), .B(n26233), .C(n30035), .D(n23537), 
         .Z(clk_enable_234)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1970_4_lut_4_lut.init = 16'hd555;
    LUT4 i1864_2_lut_2_lut (.A(resetn_c), .B(quad_set_valid_N_2333), .Z(clk_enable_315)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1864_2_lut_2_lut.init = 16'hdddd;
    LUT4 mux_158_i8_3_lut_4_lut_adj_674 (.A(n16817), .B(n30102), .C(\SLO_buf[11]_adj_312 ), 
         .D(\SLO_buf[21]_adj_313 ), .Z(\spi_data_out_r_39__N_4419[7] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i8_3_lut_4_lut_adj_674.init = 16'hf1e0;
    LUT4 i1_3_lut_4_lut_4_lut_adj_675 (.A(resetn_c), .B(EM_STOP), .C(clk_enable_256), 
         .D(n29999), .Z(clk_enable_12)) /* synthesis lut_function=((B ((D)+!C)+!B (D))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_675.init = 16'hff5d;
    LUT4 i1_4_lut_4_lut_adj_676 (.A(resetn_c), .B(n28514), .C(n23916), 
         .D(n26587), .Z(clk_enable_749)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_4_lut_adj_676.init = 16'h7555;
    LUT4 i1_4_lut_4_lut_adj_677 (.A(resetn_c), .B(n27013), .C(n23916), 
         .D(n30011), .Z(clk_enable_388)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_4_lut_adj_677.init = 16'hd555;
    LUT4 i1_2_lut_4_lut_4_lut_adj_678 (.A(resetn_c), .B(n26207), .C(n23526), 
         .D(n23916), .Z(clk_enable_898)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_4_lut_4_lut_adj_678.init = 16'hd555;
    LUT4 i1962_2_lut_4_lut_4_lut (.A(resetn_c), .B(n30062), .C(n23916), 
         .D(n26633), .Z(clk_enable_180)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1962_2_lut_4_lut_4_lut.init = 16'hd555;
    LUT4 i1_2_lut_2_lut_adj_679 (.A(resetn_c), .B(n18), .Z(n2193)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_2_lut_adj_679.init = 16'hdddd;
    LUT4 mux_158_i7_3_lut_4_lut_adj_680 (.A(n16817), .B(n30102), .C(\SLO_buf[10]_adj_314 ), 
         .D(\SLO_buf[20]_adj_315 ), .Z(\spi_data_out_r_39__N_4419[6] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i7_3_lut_4_lut_adj_680.init = 16'hf1e0;
    LUT4 i1987_4_lut_4_lut (.A(resetn_c), .B(n28540), .C(n30035), .D(n30036), 
         .Z(clk_enable_244)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1987_4_lut_4_lut.init = 16'h7555;
    LUT4 resetn_N_2923_I_0_2_lut_2_lut (.A(resetn_c), .B(clear_intrpt_adj_316), 
         .Z(intrpt_out_N_2926)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_N_2923_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_3_lut_3_lut_adj_681 (.A(resetn_c), .B(n18), .C(pwm_out_1_N_6306), 
         .Z(clk_100k_enable_1)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_3_lut_adj_681.init = 16'hfdfd;
    LUT4 reduce_or_1166_i1_4_lut_4_lut (.A(resetn_c), .B(n25889), .C(n30083), 
         .D(\quad_homing[1]_adj_317 ), .Z(n1_adj_318)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam reduce_or_1166_i1_4_lut_4_lut.init = 16'h55d5;
    LUT4 i1_2_lut_2_lut_adj_682 (.A(resetn_c), .B(n20647), .Z(clk_enable_595)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_2_lut_adj_682.init = 16'hdddd;
    LUT4 resetn_N_861_I_0_2_lut_rep_639_2_lut (.A(resetn_c), .B(EM_STOP), 
         .Z(n30039)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_N_861_I_0_2_lut_rep_639_2_lut.init = 16'hdddd;
    LUT4 mux_426_i10_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[9]), 
         .D(quad_count_adj_322[9]), .Z(\spi_data_out_r_39__N_2023[9] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_683 (.A(n30000), .B(n12), .C(\address_7__N_565[1] ), 
         .D(n28506), .Z(n25271)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_683.init = 16'h0010;
    LUT4 mux_422_i25_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[24]), 
         .D(quad_count[24]), .Z(\spi_data_out_r_39__N_1083[24] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_684 (.A(n28290), .B(n30198), .C(n32), .D(n27259), 
         .Z(clear_intrpt_N_3001)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_684.init = 16'h0100;
    LUT4 mux_426_i9_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[8]), 
         .D(quad_count_adj_322[8]), .Z(\spi_data_out_r_39__N_2023[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_422_i12_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[11]), 
         .D(quad_count[11]), .Z(\spi_data_out_r_39__N_1083[11] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_685 (.A(n30197), .B(n30196), .C(spi_cmd[0]), .D(n30195), 
         .Z(n27259)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_685.init = 16'h0200;
    LUT4 mux_426_i8_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[7]), 
         .D(quad_count_adj_322[7]), .Z(\spi_data_out_r_39__N_2023[7] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_422_i28_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[27]), 
         .D(quad_count[27]), .Z(\spi_data_out_r_39__N_1083[27] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i6_3_lut_4_lut_adj_686 (.A(n16817), .B(n30102), .C(\SLO_buf[9]_adj_275 ), 
         .D(\SLO_buf[19]_adj_282 ), .Z(\spi_data_out_r_39__N_4419[5] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i6_3_lut_4_lut_adj_686.init = 16'hf1e0;
    LUT4 mux_158_i5_3_lut_4_lut_adj_687 (.A(n16817), .B(n30102), .C(\SLO_buf[8]_adj_277 ), 
         .D(\SLO_buf[18]_adj_284 ), .Z(\spi_data_out_r_39__N_4419[4] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i5_3_lut_4_lut_adj_687.init = 16'hf1e0;
    LUT4 mux_426_i7_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[6]), 
         .D(quad_count_adj_322[6]), .Z(\spi_data_out_r_39__N_2023[6] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_701 (.A(spi_addr[2]), .B(spi_cmd[0]), .Z(n30101)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_rep_701.init = 16'heeee;
    LUT4 i1_4_lut_adj_688 (.A(n26013), .B(n26015), .C(n26007), .D(n26011), 
         .Z(n32)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_688.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut_adj_689 (.A(spi_addr[2]), .B(spi_cmd[0]), .C(spi_cmd[1]), 
         .D(spi_addr[3]), .Z(n27095)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_3_lut_4_lut_adj_689.init = 16'hfeff;
    LUT4 i1_2_lut_adj_690 (.A(spi_addr[4]), .B(spi_cmd[8]), .Z(n26013)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_adj_690.init = 16'heeee;
    LUT4 i1_2_lut_rep_702 (.A(spi_addr[1]), .B(spi_addr[0]), .Z(n30102)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_2_lut_rep_702.init = 16'hbbbb;
    LUT4 i1_3_lut_adj_691 (.A(spi_addr[5]), .B(spi_cmd[12]), .C(spi_cmd[14]), 
         .Z(n26015)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_3_lut_adj_691.init = 16'hfefe;
    LUT4 i1_2_lut_adj_692 (.A(spi_cmd[4]), .B(spi_cmd[6]), .Z(n26007)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_adj_692.init = 16'heeee;
    LUT4 i1_2_lut_adj_693 (.A(spi_cmd[13]), .B(spi_addr[6]), .Z(n26011)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_adj_693.init = 16'heeee;
    LUT4 i1_4_lut_adj_694 (.A(spi_addr[2]), .B(n24275), .C(n30156), .D(spi_cmd[0]), 
         .Z(spi_data_out_r_39__N_1868)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_4_lut_adj_694.init = 16'h1000;
    LUT4 i1_2_lut_rep_592_3_lut (.A(spi_addr[1]), .B(spi_addr[0]), .C(n16817), 
         .Z(n29992)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_2_lut_rep_592_3_lut.init = 16'hfbfb;
    LUT4 mux_158_i4_3_lut_4_lut_adj_695 (.A(n16817), .B(n30102), .C(\SLO_buf[7]_adj_279 ), 
         .D(\SLO_buf[17]_adj_286 ), .Z(\spi_data_out_r_39__N_4419[3] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i4_3_lut_4_lut_adj_695.init = 16'hf1e0;
    LUT4 mux_426_i6_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[5]), 
         .D(quad_count_adj_322[5]), .Z(\spi_data_out_r_39__N_2023[5] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_426_i25_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[24]), 
         .D(quad_count_adj_322[24]), .Z(\spi_data_out_r_39__N_2023[24] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3740_4_lut_then_4_lut (.A(spi_cmd[15]), .B(\address_7__N_549[1] ), 
         .C(n1220[9]), .D(wb_dat_o[3]), .Z(n30222)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i3740_4_lut_then_4_lut.init = 16'hfbbb;
    LUT4 mux_158_i3_3_lut_4_lut_adj_696 (.A(n16817), .B(n30102), .C(\SLO_buf[6]_adj_281 ), 
         .D(\SLO_buf[16]_adj_288 ), .Z(\spi_data_out_r_39__N_4419[2] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i3_3_lut_4_lut_adj_696.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_793 (.A(spi_cmd[11]), .B(spi_cmd[3]), .Z(n30193)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_rep_793.init = 16'heeee;
    LUT4 i1_3_lut_rep_684_4_lut (.A(spi_cmd[11]), .B(spi_cmd[3]), .C(spi_cmd[9]), 
         .D(spi_cmd[5]), .Z(n30084)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_3_lut_rep_684_4_lut.init = 16'hfffe;
    LUT4 i23750_2_lut_3_lut (.A(spi_cmd[11]), .B(spi_cmd[3]), .C(spi_cmd[1]), 
         .Z(n28452)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i23750_2_lut_3_lut.init = 16'hfefe;
    LUT4 i4_2_lut_rep_794 (.A(spi_cmd[10]), .B(spi_addr[7]), .Z(n30194)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i4_2_lut_rep_794.init = 16'heeee;
    LUT4 i1_4_lut_adj_697 (.A(n27143), .B(n30198), .C(n32), .D(n30084), 
         .Z(spi_data_out_r_39__N_5191)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_697.init = 16'h0002;
    LUT4 i1_3_lut_rep_612_4_lut (.A(spi_cmd[10]), .B(spi_addr[7]), .C(spi_cmd[7]), 
         .D(n30084), .Z(n30012)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_3_lut_rep_612_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_698 (.A(n30194), .B(spi_cmd[7]), .C(spi_addr[2]), 
         .D(n27137), .Z(n27143)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_698.init = 16'h0100;
    LUT4 i1_2_lut_rep_795 (.A(spi_cmd[15]), .B(spi_addr[2]), .Z(n30195)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_795.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_699 (.A(spi_cmd[15]), .B(spi_addr[2]), 
         .C(spi_addr[1]), .D(spi_cmd[2]), .Z(n27239)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_699.init = 16'h8000;
    LUT4 i1_2_lut_rep_796 (.A(spi_cmd[7]), .B(spi_cmd[2]), .Z(n30196)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_rep_796.init = 16'heeee;
    LUT4 i1_2_lut_rep_693_3_lut_4_lut (.A(spi_cmd[7]), .B(spi_cmd[2]), .C(spi_addr[7]), 
         .D(spi_cmd[10]), .Z(n30093)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_rep_693_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_797 (.A(spi_addr[0]), .B(spi_addr[1]), .Z(n30197)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_2_lut_rep_797.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_adj_700 (.A(spi_addr[0]), .B(spi_addr[1]), .C(spi_cmd[0]), 
         .Z(n23469)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_2_lut_3_lut_adj_700.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_701 (.A(spi_addr[0]), .B(spi_addr[1]), 
         .C(spi_addr[7]), .D(spi_cmd[10]), .Z(n27169)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_2_lut_3_lut_4_lut_adj_701.init = 16'h0002;
    LUT4 i1_2_lut_rep_798 (.A(spi_cmd[1]), .B(spi_addr[3]), .Z(n30198)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_rep_798.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut_4_lut_adj_702 (.A(spi_cmd[1]), .B(spi_addr[3]), 
         .C(spi_addr[0]), .D(spi_addr[1]), .Z(n27037)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_3_lut_4_lut_adj_702.init = 16'hffdf;
    LUT4 i1_3_lut_rep_696_4_lut (.A(spi_addr[1]), .B(spi_addr[0]), .C(spi_cmd[2]), 
         .D(spi_cmd[0]), .Z(n30096)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_3_lut_rep_696_4_lut.init = 16'hfbff;
    LUT4 i1_2_lut_rep_800 (.A(spi_addr[0]), .B(spi_addr[2]), .Z(n30200)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_2_lut_rep_800.init = 16'hbbbb;
    LUT4 i24129_4_lut (.A(n26655), .B(n30198), .C(n30154), .D(n27323), 
         .Z(spi_data_out_r_39__N_5534)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i24129_4_lut.init = 16'h0010;
    LUT4 i1_4_lut_adj_703 (.A(n30194), .B(n30084), .C(n27057), .D(spi_cmd[7]), 
         .Z(n27323)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_703.init = 16'hfffe;
    LUT4 i1_4_lut_adj_704 (.A(n28290), .B(n30198), .C(n32), .D(n27183), 
         .Z(spi_data_out_r_39__N_5877)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_704.init = 16'h0100;
    LUT4 i1_4_lut_adj_705 (.A(n30197), .B(spi_cmd[7]), .C(n27177), .D(spi_cmd[15]), 
         .Z(n27183)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_4_lut_adj_705.init = 16'h2000;
    LUT4 mux_422_i24_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[23]), 
         .D(quad_count[23]), .Z(\spi_data_out_r_39__N_1083[23] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_706 (.A(n27245), .B(n30198), .C(n32), .D(n30084), 
         .Z(spi_data_out_r_39__N_6220)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_706.init = 16'h0002;
    LUT4 i1_4_lut_adj_707 (.A(n30194), .B(spi_addr[0]), .C(spi_cmd[7]), 
         .D(n27239), .Z(n27245)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_707.init = 16'h0100;
    LUT4 mux_426_i5_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[4]), 
         .D(quad_count_adj_322[4]), .Z(\spi_data_out_r_39__N_2023[4] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_426_i24_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[23]), 
         .D(quad_count_adj_322[23]), .Z(\spi_data_out_r_39__N_2023[23] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_4_lut_adj_708 (.A(spi_cmd[15]), .B(spi_cmd[2]), .C(spi_cmd[7]), 
         .D(spi_addr[0]), .Z(n26771)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_708.init = 16'h0008;
    LUT4 mux_422_i2_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[1]), 
         .D(quad_count[1]), .Z(\spi_data_out_r_39__N_1083[1] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_811 (.A(mem_burst_cnt[1]), .B(mem_burst_cnt[4]), .Z(n30211)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(355[47:82])
    defparam i1_2_lut_rep_811.init = 16'heeee;
    LUT4 i1_3_lut_rep_692_4_lut (.A(mem_burst_cnt[1]), .B(mem_burst_cnt[4]), 
         .C(n18233), .D(n23343), .Z(n30092)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/s_links/sources/spi_ctrl.v(355[47:82])
    defparam i1_3_lut_rep_692_4_lut.init = 16'hffef;
    LUT4 i5903_2_lut_rep_812 (.A(spi_cmd[15]), .B(\address_7__N_549[1] ), 
         .Z(n30212)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i5903_2_lut_rep_812.init = 16'h4444;
    LUT4 i346_2_lut_3_lut (.A(spi_cmd[15]), .B(\address_7__N_549[1] ), .C(spi_addr_valid_N_732), 
         .Z(n1277)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i346_2_lut_3_lut.init = 16'h4040;
    LUT4 i24101_2_lut_3_lut (.A(spi_cmd[15]), .B(\address_7__N_549[1] ), 
         .C(n1220[10]), .Z(n11068)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i24101_2_lut_3_lut.init = 16'hbfbf;
    LUT4 mux_422_i27_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[26]), 
         .D(quad_count[26]), .Z(\spi_data_out_r_39__N_1083[26] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_709 (.A(n26257), .B(n23469), .C(n24312), .D(n29997), 
         .Z(spi_data_out_r_39__N_1398)) /* synthesis lut_function=(!(A ((C)+!B)+!A ((C (D))+!B))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_4_lut_adj_709.init = 16'h0c4c;
    LUT4 mux_422_i26_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[25]), 
         .D(quad_count[25]), .Z(\spi_data_out_r_39__N_1083[25] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_422_i31_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[30]), 
         .D(quad_count[30]), .Z(\spi_data_out_r_39__N_1083[30] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut_adj_710 (.A(n30013), .B(n30198), .C(n26641), .D(n30084), 
         .Z(n24312)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_710.init = 16'hfffe;
    LUT4 mux_426_i4_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[3]), 
         .D(quad_count_adj_322[3]), .Z(\spi_data_out_r_39__N_2023[3] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_158_i2_3_lut_4_lut_adj_711 (.A(n16817), .B(n30102), .C(\SLO_buf[5]_adj_319 ), 
         .D(\SLO_buf[15]_adj_290 ), .Z(\spi_data_out_r_39__N_4419[1] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_158_i2_3_lut_4_lut_adj_711.init = 16'hf1e0;
    FD1P3IX spi_byte_cnt_1788__i2 (.D(n21[2]), .SP(clk_enable_915), .CD(n12446), 
            .CK(clk), .Q(spi_byte_cnt[2]));   // c:/s_links/sources/spi_ctrl.v(383[46:62])
    defparam spi_byte_cnt_1788__i2.GSR = "ENABLED";
    FD1P3IX spi_byte_cnt_1788__i3 (.D(n21[3]), .SP(clk_enable_915), .CD(n12446), 
            .CK(clk), .Q(spi_byte_cnt[3]));   // c:/s_links/sources/spi_ctrl.v(383[46:62])
    defparam spi_byte_cnt_1788__i3.GSR = "ENABLED";
    LUT4 mux_426_i3_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[2]), 
         .D(quad_count_adj_322[2]), .Z(\spi_data_out_r_39__N_2023[2] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 wb_xfer_done_I_0_238_2_lut_rep_816 (.A(\address_7__N_549[1] ), .B(wb_dat_o[4]), 
         .Z(n30216)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_ctrl.v(347[31:57])
    defparam wb_xfer_done_I_0_238_2_lut_rep_816.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_712 (.A(\address_7__N_549[1] ), .B(wb_dat_o[4]), 
         .C(n1220[11]), .D(spi_cmd[15]), .Z(clk_enable_756)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(347[31:57])
    defparam i1_2_lut_3_lut_4_lut_adj_712.init = 16'h8000;
    LUT4 i1_3_lut_4_lut_4_lut_adj_713 (.A(\address_7__N_549[1] ), .B(wb_dat_o[4]), 
         .C(n1220[3]), .D(n30059), .Z(n24466)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(347[31:57])
    defparam i1_3_lut_4_lut_4_lut_adj_713.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_adj_714 (.A(\address_7__N_549[1] ), .B(wb_dat_o[4]), 
         .C(spi_idle), .Z(n26661)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(347[31:57])
    defparam i1_2_lut_3_lut_adj_714.init = 16'h0808;
    PFUMX i59 (.BLUT(n24197), .ALUT(rd_en_N_717), .C0(n1220[9]), .Z(n26));
    LUT4 i1_2_lut_3_lut_adj_715 (.A(\address_7__N_549[1] ), .B(wb_dat_o[4]), 
         .C(n1220[11]), .Z(n6)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(347[31:57])
    defparam i1_2_lut_3_lut_adj_715.init = 16'h7070;
    FD1P3IX spi_byte_cnt_1788__i1 (.D(n21[1]), .SP(clk_enable_915), .CD(n12446), 
            .CK(clk), .Q(spi_byte_cnt[1]));   // c:/s_links/sources/spi_ctrl.v(383[46:62])
    defparam spi_byte_cnt_1788__i1.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_716 (.A(\address_7__N_549[1] ), .B(wb_dat_o[4]), 
         .C(n1220[10]), .D(spi_cmd[15]), .Z(n26715)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(347[31:57])
    defparam i1_2_lut_3_lut_4_lut_adj_716.init = 16'h0800;
    LUT4 i13340_2_lut_3_lut_3_lut (.A(\address_7__N_549[1] ), .B(wb_dat_o[4]), 
         .C(n30059), .Z(wr_en_N_701)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(347[31:57])
    defparam i13340_2_lut_3_lut_3_lut.init = 16'h0808;
    LUT4 mux_426_i2_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[1]), 
         .D(quad_count_adj_322[1]), .Z(\spi_data_out_r_39__N_2023[1] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_597_4_lut (.A(n30194), .B(n30084), .C(spi_cmd[7]), 
         .D(n30013), .Z(n29997)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_rep_597_4_lut.init = 16'hfffe;
    LUT4 mux_422_i11_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[10]), 
         .D(quad_count[10]), .Z(\spi_data_out_r_39__N_1083[10] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 wb_xfer_done_I_0_242_2_lut_rep_817 (.A(\address_7__N_549[1] ), .B(wb_dat_o[3]), 
         .Z(n30217)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_ctrl.v(288[31:57])
    defparam wb_xfer_done_I_0_242_2_lut_rep_817.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_717 (.A(\address_7__N_549[1] ), .B(wb_dat_o[3]), 
         .C(n1220[7]), .Z(n26765)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(288[31:57])
    defparam i1_2_lut_3_lut_adj_717.init = 16'h8080;
    LUT4 i1_2_lut_rep_613 (.A(spi_cmd[15]), .B(n32), .Z(n30013)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_rep_613.init = 16'hdddd;
    LUT4 spi_xfer_done_bdd_3_lut_3_lut (.A(\address_7__N_549[1] ), .B(wb_dat_o[3]), 
         .C(wb_dat_o[4]), .Z(n29911)) /* synthesis lut_function=(A (B+!(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(288[31:57])
    defparam spi_xfer_done_bdd_3_lut_3_lut.init = 16'h8a8a;
    LUT4 i3641_4_lut_4_lut (.A(\address_7__N_549[1] ), .B(wb_dat_o[3]), 
         .C(n1220[3]), .D(n1220[4]), .Z(n7963)) /* synthesis lut_function=(A (B (C))+!A (D)) */ ;   // c:/s_links/sources/spi_ctrl.v(288[31:57])
    defparam i3641_4_lut_4_lut.init = 16'hd580;
    LUT4 spi_xfer_done_bdd_2_lut_24373_3_lut (.A(\address_7__N_549[1] ), .B(wb_dat_o[3]), 
         .C(n1220[7]), .Z(n29910)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(288[31:57])
    defparam spi_xfer_done_bdd_2_lut_24373_3_lut.init = 16'h0808;
    LUT4 mux_426_i1_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[0]), 
         .D(quad_count_adj_322[0]), .Z(\spi_data_out_r_39__N_2023[0] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_426_i23_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[22]), 
         .D(quad_count_adj_322[22]), .Z(\spi_data_out_r_39__N_2023[22] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3695_2_lut_3_lut (.A(\address_7__N_549[1] ), .B(n30059), .C(n1220[9]), 
         .Z(n8019)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i3695_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_4_lut_adj_718 (.A(clk_enable_627), .B(EM_STOP), .C(n30007), 
         .D(n30016), .Z(clk_enable_38)) /* synthesis lut_function=(A+!((C (D))+!B)) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_adj_718.init = 16'haeee;
    LUT4 i23917_3_lut (.A(n25271), .B(n4382), .C(n28534), .Z(n5327[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i23917_3_lut.init = 16'hcaca;
    LUT4 mux_426_i22_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[21]), 
         .D(quad_count_adj_322[21]), .Z(\spi_data_out_r_39__N_2023[21] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_620 (.A(resetn_c), .B(n18654), .Z(n30020)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/mcm_top.v(17[27:33])
    defparam i1_2_lut_rep_620.init = 16'h8888;
    LUT4 mux_426_i32_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[31]), 
         .D(quad_count_adj_322[31]), .Z(\spi_data_out_r_39__N_2023[31] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i16352_1_lut_2_lut (.A(resetn_c), .B(n18654), .Z(clk_enable_227)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/s_links/sources/mcm_top.v(17[27:33])
    defparam i16352_1_lut_2_lut.init = 16'h7777;
    LUT4 mux_426_i31_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[30]), 
         .D(quad_count_adj_322[30]), .Z(\spi_data_out_r_39__N_2023[30] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3676_4_lut (.A(mem_rdata_update_N_729), .B(n30074), .C(\address_7__N_549[1] ), 
         .D(clk_enable_756), .Z(n8000)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i3676_4_lut.init = 16'h3b0a;
    LUT4 i1_2_lut_3_lut_4_lut_adj_719 (.A(\address_7__N_549[1] ), .B(n23860), 
         .C(n28506), .D(n30136), .Z(n25421)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C+(D))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_719.init = 16'hf7f0;
    LUT4 mux_426_i30_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[29]), 
         .D(quad_count_adj_322[29]), .Z(\spi_data_out_r_39__N_2023[29] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_422_i29_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[28]), 
         .D(quad_count[28]), .Z(\spi_data_out_r_39__N_1083[28] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3635_4_lut_4_lut (.A(\address_7__N_549[1] ), .B(n23860), .C(n1220[6]), 
         .D(n1220[7]), .Z(n7957)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (D)) */ ;
    defparam i3635_4_lut_4_lut.init = 16'hf7a0;
    LUT4 i1_4_lut_adj_720 (.A(n1220[11]), .B(n11727), .C(n26333), .D(n7970), 
         .Z(n11728)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_720.init = 16'hecee;
    LUT4 i1_4_lut_adj_721 (.A(\address_7__N_549[1] ), .B(spi_cmd[15]), .C(mem_rdata_update_N_729), 
         .D(spi_addr_valid_N_732), .Z(n11727)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_721.init = 16'ha8a0;
    LUT4 i1_4_lut_adj_722 (.A(spi_cmd[15]), .B(\address_7__N_549[1] ), .C(n30169), 
         .D(n26661), .Z(n26333)) /* synthesis lut_function=(!(A (B)+!A (B (C+!(D))))) */ ;
    defparam i1_4_lut_adj_722.init = 16'h3733;
    LUT4 i3643_4_lut_4_lut (.A(\address_7__N_549[1] ), .B(n23860), .C(n1220[2]), 
         .D(n1220[3]), .Z(n7965)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (D)) */ ;
    defparam i3643_4_lut_4_lut.init = 16'hf7a0;
    LUT4 i1_4_lut_adj_723 (.A(n30060), .B(n25457), .C(\address_7__N_549[1] ), 
         .D(n24198), .Z(n24197)) /* synthesis lut_function=(!(A+!(B (C)+!B !((D)+!C)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_723.init = 16'h4050;
    LUT4 i1_4_lut_adj_724 (.A(n30074), .B(n8019), .C(n1277), .D(n11068), 
         .Z(n24505)) /* synthesis lut_function=(A (B+(C))+!A (B+(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_724.init = 16'hfcfd;
    LUT4 i3629_4_lut (.A(spi_addr_valid_N_732), .B(n26765), .C(\address_7__N_549[1] ), 
         .D(n30074), .Z(n7951)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A ((D)+!B))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i3629_4_lut.init = 16'h0ace;
    LUT4 i1_4_lut_adj_725 (.A(n26043), .B(n1220[7]), .C(n30017), .D(n30216), 
         .Z(n24758)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_725.init = 16'heaaa;
    LUT4 i1_4_lut_adj_726 (.A(spi_cmd_cnt), .B(n1220[6]), .C(n23412), 
         .D(\address_7__N_549[1] ), .Z(n26043)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_726.init = 16'ha0ec;
    LUT4 i1_4_lut_adj_727 (.A(spi_cmd_cnt), .B(n24466), .C(n8), .D(n23412), 
         .Z(n24465)) /* synthesis lut_function=(A (B+(C))+!A (B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_727.init = 16'hfdfc;
    LUT4 i1_2_lut_3_lut_adj_728 (.A(spi_cmd[0]), .B(n30084), .C(spi_cmd[15]), 
         .Z(n26467)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_3_lut_adj_728.init = 16'hdfdf;
    LUT4 i1_4_lut_adj_729 (.A(n30012), .B(n30198), .C(n26655), .D(spi_cmd[15]), 
         .Z(n26483)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_4_lut_adj_729.init = 16'hfeff;
    LUT4 i1_2_lut_4_lut_adj_730 (.A(n30194), .B(n30084), .C(n30161), .D(spi_cmd[15]), 
         .Z(n26599)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_4_lut_adj_730.init = 16'hfeff;
    LUT4 mux_426_i29_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[28]), 
         .D(quad_count_adj_322[28]), .Z(\spi_data_out_r_39__N_2023[28] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_adj_731 (.A(spi_addr[2]), .B(n32), .Z(n26655)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_adj_731.init = 16'hdddd;
    LUT4 i14_3_lut (.A(n1220[2]), .B(spi_cmd_start_reg_N_746), .C(\address_7__N_549[1] ), 
         .Z(n8)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i14_3_lut.init = 16'hcaca;
    LUT4 i3653_4_lut (.A(spi_cmd_start_reg_N_746), .B(\address_7__N_565[1] ), 
         .C(\address_7__N_549[1] ), .D(spi_cmd_start_reg_N_745), .Z(n7977)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i3653_4_lut.init = 16'hce0a;
    LUT4 mux_426_i28_3_lut_4_lut (.A(n30200), .B(n23623), .C(quad_buffer_adj_321[27]), 
         .D(quad_count_adj_322[27]), .Z(\spi_data_out_r_39__N_2023[27] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_426_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_422_i22_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[21]), 
         .D(quad_count[21]), .Z(\spi_data_out_r_39__N_1083[21] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n22554_bdd_4_lut_24464 (.A(n22554), .B(pwm), .C(n4_adj_320), 
         .D(\status_cntr[11] ), .Z(n29985)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam n22554_bdd_4_lut_24464.init = 16'hf0ee;
    LUT4 i15_4_lut (.A(n1220[11]), .B(\address_7__N_549[1] ), .C(spi_addr_valid_N_732), 
         .D(n30113), .Z(clk_enable_321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i15_4_lut.init = 16'hcfca;
    LUT4 mux_422_i1_3_lut_4_lut (.A(n23623), .B(n30159), .C(quad_buffer[0]), 
         .D(quad_count[0]), .Z(\spi_data_out_r_39__N_1083[0] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_422_i1_3_lut_4_lut.init = 16'hf1e0;
    FD1P3IX mem_burst_cnt_1790__i2 (.D(n37_adj_7039[2]), .SP(clk_enable_1128), 
            .CD(n12460), .CK(clk), .Q(mem_burst_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_1790__i2.GSR = "ENABLED";
    FD1P3IX mem_burst_cnt_1790__i7 (.D(n37_adj_7039[7]), .SP(clk_enable_1128), 
            .CD(n12460), .CK(clk), .Q(mem_burst_cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_1790__i7.GSR = "ENABLED";
    FD1P3IX mem_burst_cnt_1790__i1 (.D(n37_adj_7039[1]), .SP(clk_enable_1128), 
            .CD(n12460), .CK(clk), .Q(mem_burst_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_1790__i1.GSR = "ENABLED";
    FD1P3IX mem_burst_cnt_1790__i6 (.D(n37_adj_7039[6]), .SP(clk_enable_1128), 
            .CD(n12460), .CK(clk), .Q(mem_burst_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_1790__i6.GSR = "ENABLED";
    FD1P3IX mem_burst_cnt_1790__i5 (.D(n37_adj_7039[5]), .SP(clk_enable_1128), 
            .CD(n12460), .CK(clk), .Q(mem_burst_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_1790__i5.GSR = "ENABLED";
    FD1P3IX mem_burst_cnt_1790__i4 (.D(n37_adj_7039[4]), .SP(clk_enable_1128), 
            .CD(n12460), .CK(clk), .Q(mem_burst_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_1790__i4.GSR = "ENABLED";
    FD1P3IX mem_burst_cnt_1790__i3 (.D(n37_adj_7039[3]), .SP(clk_enable_1128), 
            .CD(n12460), .CK(clk), .Q(mem_burst_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_1790__i3.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_713 (.A(spi_cmd_start_reg_N_745), .B(n1220[9]), .Z(n30113)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_713.init = 16'heeee;
    LUT4 i11_3_lut_4_lut (.A(spi_cmd_start_reg_N_745), .B(n1220[9]), .C(n1220[10]), 
         .D(n30212), .Z(clk_enable_1110)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam i11_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i13909_2_lut_3_lut (.A(spi_cmd_start_reg_N_745), .B(n1220[9]), 
         .C(n1220[10]), .Z(n18232)) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;
    defparam i13909_2_lut_3_lut.init = 16'h0e0e;
    FD1P3IX spi_cmd_valid_223 (.D(spi_cmd_cnt), .SP(clk_enable_1106), .CD(n18231), 
            .CK(clk), .Q(spi_cmd_valid)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_valid_223.GSR = "ENABLED";
    FD1P3IX spi_data_valid_226 (.D(spi_data_valid_N_737), .SP(clk_enable_1110), 
            .CD(n18232), .CK(clk), .Q(spi_data_valid)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data_valid_226.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut_adj_732 (.A(spi_cmd[15]), .B(spi_byte_cnt[3]), .C(n27365), 
         .D(n30127), .Z(clk_enable_569)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_4_lut_adj_732.init = 16'h1000;
    LUT4 i334_2_lut_rep_723 (.A(\address_7__N_549[1] ), .B(n1220[4]), .Z(n30123)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i334_2_lut_rep_723.init = 16'h8888;
    LUT4 i23972_2_lut_3_lut (.A(\address_7__N_549[1] ), .B(n1220[4]), .C(spi_cmd_cnt), 
         .Z(clk_enable_867)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i23972_2_lut_3_lut.init = 16'h0808;
    LUT4 i4311_2_lut_3_lut (.A(\address_7__N_549[1] ), .B(n1220[4]), .C(spi_cmd_cnt), 
         .Z(clk_enable_859)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i4311_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_3_lut_4_lut_adj_733 (.A(spi_cmd[2]), .B(spi_addr[1]), .C(spi_cmd[15]), 
         .D(spi_addr[0]), .Z(n27223)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut_adj_733.init = 16'h0080;
    LUT4 i1477_3_lut_rep_727 (.A(spi_cmd_start_reg_N_745), .B(\address_7__N_549[1] ), 
         .C(n1220[10]), .Z(n30127)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1477_3_lut_rep_727.init = 16'hcaca;
    LUT4 i1_2_lut_rep_654_4_lut (.A(spi_cmd_start_reg_N_745), .B(\address_7__N_549[1] ), 
         .C(n1220[10]), .D(spi_cmd[15]), .Z(n30054)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_2_lut_rep_654_4_lut.init = 16'h00ca;
    FD1P3IX mem_burst_cnt_1790__i0 (.D(n37_adj_7039[0]), .SP(clk_enable_1128), 
            .CD(n12460), .CK(clk), .Q(mem_burst_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_1790__i0.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_735 (.A(n1220[5]), .B(spi_cmd_start_reg_N_746), .Z(n30135)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_2_lut_rep_735.init = 16'heeee;
    LUT4 i1_2_lut_rep_660_3_lut (.A(n1220[5]), .B(spi_cmd_start_reg_N_746), 
         .C(n1220[4]), .Z(n30060)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_2_lut_rep_660_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_736 (.A(n1220[7]), .B(n1220[3]), .Z(n30136)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_2_lut_rep_736.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_734 (.A(n1220[7]), .B(n1220[3]), .C(n1220[9]), 
         .D(n30217), .Z(n4382)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_3_lut_4_lut_adj_734.init = 16'hfe00;
    LUT4 i2_2_lut_rep_600_3_lut_4_lut (.A(n1220[7]), .B(n1220[3]), .C(n23860), 
         .D(\address_7__N_549[1] ), .Z(n30000)) /* synthesis lut_function=(!(A (C (D))+!A ((C (D))+!B))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i2_2_lut_rep_600_3_lut_4_lut.init = 16'h0eee;
    LUT4 i2_2_lut_3_lut (.A(n1220[7]), .B(n1220[3]), .C(n23860), .Z(n10254)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i2_2_lut_3_lut.init = 16'he0e0;
    LUT4 i23804_2_lut_3_lut (.A(n1220[2]), .B(n1220[6]), .C(mem_rdata_update_N_729), 
         .Z(n28506)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i23804_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_3_lut_4_lut_adj_735 (.A(n1220[2]), .B(n1220[6]), .C(mem_rdata_update_N_729), 
         .D(spi_addr_valid_N_732), .Z(n25457)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_3_lut_4_lut_adj_735.init = 16'hfffe;
    LUT4 i3823_4_lut_4_lut (.A(n1220[10]), .B(\address_7__N_549[1] ), .C(n11759), 
         .D(spi_cmd[15]), .Z(address_7__N_359[0])) /* synthesis lut_function=(A ((D)+!B)+!A !(B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i3823_4_lut_4_lut.init = 16'hbf37;
    LUT4 i24159_2_lut_3_lut (.A(n1220[10]), .B(\address_7__N_549[1] ), .C(n11759), 
         .Z(n28577)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i24159_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i5068_3_lut_3_lut_3_lut (.A(n1220[10]), .B(\address_7__N_549[1] ), 
         .C(spi_cmd[15]), .Z(n9392)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i5068_3_lut_3_lut_3_lut.init = 16'h4c4c;
    LUT4 i11_3_lut_4_lut_adj_736 (.A(spi_cmd_start_reg_N_745), .B(n1220[5]), 
         .C(n1220[4]), .D(\address_7__N_549[1] ), .Z(clk_enable_1106)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam i11_3_lut_4_lut_adj_736.init = 16'hfe0e;
    LUT4 i13908_2_lut_3_lut (.A(spi_cmd_start_reg_N_745), .B(n1220[5]), 
         .C(n1220[4]), .Z(n18231)) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;
    defparam i13908_2_lut_3_lut.init = 16'h0e0e;
    LUT4 i1_2_lut_rep_745 (.A(spi_cmd[7]), .B(spi_cmd[0]), .Z(n30145)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_rep_745.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_737 (.A(spi_cmd[7]), .B(spi_cmd[0]), .C(n30084), 
         .D(n30194), .Z(n27027)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_3_lut_4_lut_adj_737.init = 16'hfffe;
    LUT4 i17490_2_lut_3_lut (.A(spi_byte_cnt[1]), .B(spi_byte_cnt[0]), .C(spi_byte_cnt[2]), 
         .Z(n21[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(383[46:62])
    defparam i17490_2_lut_3_lut.init = 16'h7878;
    LUT4 i17497_3_lut_4_lut (.A(spi_byte_cnt[1]), .B(spi_byte_cnt[0]), .C(spi_byte_cnt[2]), 
         .D(spi_byte_cnt[3]), .Z(n21[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/s_links/sources/spi_ctrl.v(383[46:62])
    defparam i17497_3_lut_4_lut.init = 16'h7f80;
    LUT4 i1_2_lut_rep_747 (.A(spi_cmd[0]), .B(spi_addr[1]), .Z(n30147)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_2_lut_rep_747.init = 16'h2222;
    LUT4 i1_3_lut_4_lut_adj_738 (.A(spi_cmd[0]), .B(spi_addr[1]), .C(n24275), 
         .D(n30200), .Z(spi_data_out_r_39__N_2103)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_3_lut_4_lut_adj_738.init = 16'h0002;
    LUT4 i1_3_lut_4_lut_adj_739 (.A(spi_cmd[0]), .B(spi_addr[1]), .C(n30159), 
         .D(n24275), .Z(spi_data_out_r_39__N_1163)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_3_lut_4_lut_adj_739.init = 16'h0002;
    LUT4 mux_428_i1_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[0]), 
         .D(quad_count_adj_324[0]), .Z(\spi_data_out_r_39__N_2493[0] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i32_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[31]), 
         .D(quad_count_adj_324[31]), .Z(\spi_data_out_r_39__N_2493[31] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_428_i31_3_lut_4_lut (.A(n16815), .B(n30200), .C(quad_buffer_adj_323[30]), 
         .D(quad_count_adj_324[30]), .Z(\spi_data_out_r_39__N_2493[30] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mux_428_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_4_lut_adj_740 (.A(spi_addr[3]), .B(spi_cmd[1]), .C(spi_cmd[2]), 
         .D(spi_addr[2]), .Z(n26263)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_3_lut_4_lut_adj_740.init = 16'hefff;
    LUT4 i1_3_lut_4_lut_adj_741 (.A(spi_addr[3]), .B(spi_cmd[1]), .C(spi_addr[2]), 
         .D(spi_cmd[2]), .Z(n26257)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_3_lut_4_lut_adj_741.init = 16'hfeff;
    LUT4 i1_3_lut_4_lut_adj_742 (.A(spi_cmd[0]), .B(spi_addr[1]), .C(n24275), 
         .D(n30159), .Z(spi_data_out_r_39__N_1633)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_3_lut_4_lut_adj_742.init = 16'h0008;
    LUT4 i1_3_lut_4_lut_adj_743 (.A(spi_cmd[0]), .B(spi_addr[1]), .C(n24275), 
         .D(n30200), .Z(spi_data_out_r_39__N_2573)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_3_lut_4_lut_adj_743.init = 16'h0008;
    PFUMX i24397 (.BLUT(n30224), .ALUT(n30225), .C0(spi_cmd_start_reg_N_746), 
          .Z(n30226));
    LUT4 i1_2_lut_rep_754 (.A(spi_cmd[15]), .B(spi_cmd[2]), .Z(n30154)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_754.init = 16'h8888;
    PFUMX i24395 (.BLUT(n30221), .ALUT(n30222), .C0(n1220[10]), .Z(n30223));
    
endmodule
//
// Verilog Description of module \stepper(DEV_ID=1,UART_ADDRESS_WIDTH=4) 
//

module \stepper(DEV_ID=1,UART_ADDRESS_WIDTH=4)  (reset_r, clk, clk_enable_12, 
            n30185, n29999, clk_1MHz, GND_net, resetn_c, pin_io_c_18, 
            n30098, spi_data_out_r_39__N_4168, \spi_data_out_r_39__N_4419[0] , 
            clk_enable_759, \spi_data_r[0] , \SLO_buf[0] , n29992, \SLO_buf[13] , 
            \SLO_buf[12] , \SLO_buf[11] , \SLO_buf[10] , \spi_data_out_r_39__N_4419[35] , 
            \spi_data_out_r_39__N_4419[34] , \spi_data_out_r_39__N_4419[33] , 
            \spi_data_out_r_39__N_4419[32] , \spi_data_out_r_39__N_4419[15] , 
            \spi_data_out_r_39__N_4419[14] , \spi_data_out_r_39__N_4419[13] , 
            \spi_data_out_r_39__N_4419[12] , \spi_data_out_r_39__N_4419[11] , 
            \spi_data_out_r_39__N_4419[10] , \spi_data_out_r_39__N_4419[9] , 
            \spi_data_out_r_39__N_4419[8] , \spi_data_out_r_39__N_4419[7] , 
            \spi_data_out_r_39__N_4419[6] , \spi_data_out_r_39__N_4419[5] , 
            \spi_data_out_r_39__N_4419[4] , \spi_data_out_r_39__N_4419[3] , 
            \spi_data_out_r_39__N_4419[2] , \spi_data_out_r_39__N_4419[1] , 
            \quad_homing[0] , pin_io_c_14, n25877, spi_data_out_r_39__N_4208, 
            spi_data_out_r_39__N_4505, digital_output_r, clk_enable_256, 
            n28555, \quad_a[1] , pin_io_out_19, \quad_b[1] , uart_slot_en, 
            n30095, n28, \spi_data_r[1] , \spi_data_r[2] , \SLO_buf[1] , 
            \SLO_buf[2] , \SLO_buf[3] , \SLO_buf[4] , \SLO_buf[5] , 
            \SLO_buf[6] , \SLO_buf[7] , \SLO_buf[8] , \SLO_buf[9] , 
            \SLO_buf[14] , \SLO_buf[15] , \SLO_buf[16] , \SLO_buf[17] , 
            \SLO_buf[18] , \SLO_buf[19] , \SLO_buf[20] , \SLO_buf[21] , 
            \SLO_buf[22] , \SLO_buf[23] , \SLO_buf[24] , \SLO_buf[25] , 
            \SLO_buf[26] , \SLO_buf[27] , \SLO_buf[28] , \SLO_buf[29] , 
            NSL, UC_TXD0_c, OW_ID_N_4461, OW_ID_N_4467, n30050, n30041, 
            n30075, pin_io_c_13, \pin_intrpt[4] , pin_io_out_15, n29944, 
            pin_io_c_12, \pin_intrpt[3] , \pin_intrpt[5] , n7277, ENC_O_N_4469, 
            n30118, n30049, \mode[2] , n9) /* synthesis syn_module_defined=1 */ ;
    output reset_r;
    input clk;
    input clk_enable_12;
    input n30185;
    input n29999;
    input clk_1MHz;
    input GND_net;
    input resetn_c;
    input pin_io_c_18;
    output n30098;
    output [39:0]spi_data_out_r_39__N_4168;
    input \spi_data_out_r_39__N_4419[0] ;
    input clk_enable_759;
    input \spi_data_r[0] ;
    output \SLO_buf[0] ;
    input n29992;
    output \SLO_buf[13] ;
    output \SLO_buf[12] ;
    output \SLO_buf[11] ;
    output \SLO_buf[10] ;
    input \spi_data_out_r_39__N_4419[35] ;
    input \spi_data_out_r_39__N_4419[34] ;
    input \spi_data_out_r_39__N_4419[33] ;
    input \spi_data_out_r_39__N_4419[32] ;
    input \spi_data_out_r_39__N_4419[15] ;
    input \spi_data_out_r_39__N_4419[14] ;
    input \spi_data_out_r_39__N_4419[13] ;
    input \spi_data_out_r_39__N_4419[12] ;
    input \spi_data_out_r_39__N_4419[11] ;
    input \spi_data_out_r_39__N_4419[10] ;
    input \spi_data_out_r_39__N_4419[9] ;
    input \spi_data_out_r_39__N_4419[8] ;
    input \spi_data_out_r_39__N_4419[7] ;
    input \spi_data_out_r_39__N_4419[6] ;
    input \spi_data_out_r_39__N_4419[5] ;
    input \spi_data_out_r_39__N_4419[4] ;
    input \spi_data_out_r_39__N_4419[3] ;
    input \spi_data_out_r_39__N_4419[2] ;
    input \spi_data_out_r_39__N_4419[1] ;
    input \quad_homing[0] ;
    input pin_io_c_14;
    output n25877;
    output spi_data_out_r_39__N_4208;
    input spi_data_out_r_39__N_4505;
    output digital_output_r;
    input clk_enable_256;
    input n28555;
    output \quad_a[1] ;
    input pin_io_out_19;
    output \quad_b[1] ;
    input [3:0]uart_slot_en;
    input n30095;
    output n28;
    input \spi_data_r[1] ;
    input \spi_data_r[2] ;
    output \SLO_buf[1] ;
    output \SLO_buf[2] ;
    output \SLO_buf[3] ;
    output \SLO_buf[4] ;
    output \SLO_buf[5] ;
    output \SLO_buf[6] ;
    output \SLO_buf[7] ;
    output \SLO_buf[8] ;
    output \SLO_buf[9] ;
    output \SLO_buf[14] ;
    output \SLO_buf[15] ;
    output \SLO_buf[16] ;
    output \SLO_buf[17] ;
    output \SLO_buf[18] ;
    output \SLO_buf[19] ;
    output \SLO_buf[20] ;
    output \SLO_buf[21] ;
    output \SLO_buf[22] ;
    output \SLO_buf[23] ;
    output \SLO_buf[24] ;
    output \SLO_buf[25] ;
    output \SLO_buf[26] ;
    output \SLO_buf[27] ;
    output \SLO_buf[28] ;
    output \SLO_buf[29] ;
    output NSL;
    input UC_TXD0_c;
    output OW_ID_N_4461;
    output OW_ID_N_4467;
    output n30050;
    output n30041;
    output n30075;
    input pin_io_c_13;
    output \pin_intrpt[4] ;
    input pin_io_out_15;
    output n29944;
    input pin_io_c_12;
    output \pin_intrpt[3] ;
    output \pin_intrpt[5] ;
    output n7277;
    output ENC_O_N_4469;
    output n30118;
    output n30049;
    input \mode[2] ;
    output n9;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire clk_1MHz /* synthesis SET_AS_NETWORK=clk_1MHz, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(136[6:14])
    wire \pin_intrpt[5]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[5] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    wire [7:0]Cnt;   // c:/s_links/sources/slot_cards/stepper.v(62[11:14])
    
    wire clk_1MHz_enable_41;
    wire [7:0]n199;
    wire [51:0]SLO;   // c:/s_links/sources/slot_cards/stepper.v(63[12:15])
    
    wire clk_enable_1120, n12287, n18662, n18586;
    wire [31:0]n153;
    
    wire n11629, n30034, n10368;
    wire [11:0]n93;
    wire [11:0]n53;
    wire [11:0]Cnt_NSL;   // c:/s_links/sources/slot_cards/stepper.v(61[12:19])
    
    wire prev_MA_Temp, MA_Temp, prev_MA;
    wire [2:0]mode;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    wire n30103, n26373, n30038, n30108, n30107, clk_1MHz_enable_70, 
        n29611, SLO_buf_51__N_4358, n29610;
    wire [51:0]SLO_buf;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire clk_1MHz_enable_42, MA_Temp_N_4487, n30042, NSL_N_4500, OW_ID_N_4462, 
        n10_adj_6707, n21927, n26297, n21926, n30104, n30105, n30106, 
        n18478, n21925, n21924, n21923, n21922, n21921, n21920, 
        n21919, n21918, n25214, n24765;
    
    FD1P3IX reset_r_491 (.D(n29999), .SP(clk_enable_12), .CD(n30185), 
            .CK(clk), .Q(reset_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam reset_r_491.GSR = "DISABLED";
    FD1P3IX Cnt__i0 (.D(n199[0]), .SP(clk_1MHz_enable_41), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i0.GSR = "DISABLED";
    FD1P3IX SLO__i12 (.D(SLO[10]), .SP(clk_enable_1120), .CD(GND_net), 
            .CK(clk), .Q(SLO[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i12.GSR = "DISABLED";
    FD1P3IX SLO__i45 (.D(SLO[43]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i45.GSR = "DISABLED";
    FD1P3IX SLO__i46 (.D(SLO[44]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i46.GSR = "DISABLED";
    FD1P3IX SLO__i31 (.D(SLO[29]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i31.GSR = "DISABLED";
    LUT4 i13249_2_lut_3_lut (.A(n18662), .B(n18586), .C(n153[4]), .Z(n199[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13249_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_3_lut_rep_634 (.A(Cnt[4]), .B(n11629), .C(Cnt[1]), .Z(n30034)) /* synthesis lut_function=((B+!(C))+!A) */ ;
    defparam i1_3_lut_rep_634.init = 16'hdfdf;
    FD1P3IX SLO__i13 (.D(SLO[11]), .SP(clk_enable_1120), .CD(GND_net), 
            .CK(clk), .Q(SLO[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i13.GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut (.A(Cnt[4]), .B(n11629), .C(Cnt[1]), .D(Cnt[5]), 
         .Z(n10368)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i1_2_lut_4_lut.init = 16'hffdf;
    FD1P3IX SLO__i32 (.D(SLO[30]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i32.GSR = "DISABLED";
    FD1P3IX SLO__i33 (.D(SLO[31]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i33.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1779__i0 (.D(n53[0]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779__i0.GSR = "DISABLED";
    FD1P3IX SLO__i14 (.D(SLO[12]), .SP(clk_enable_1120), .CD(GND_net), 
            .CK(clk), .Q(SLO[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i14.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1779__i11 (.D(n53[11]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779__i11.GSR = "DISABLED";
    FD1P3IX SLO__i34 (.D(SLO[32]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i34.GSR = "DISABLED";
    FD1P3IX SLO__i35 (.D(SLO[33]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i35.GSR = "DISABLED";
    FD1P3IX SLO__i1 (.D(pin_io_c_18), .SP(clk_enable_1120), .CD(GND_net), 
            .CK(clk), .Q(SLO[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i1.GSR = "DISABLED";
    FD1P3IX SLO__i44 (.D(SLO[42]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i44.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1779__i10 (.D(n53[10]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779__i10.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1779__i9 (.D(n53[9]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779__i9.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1779__i8 (.D(n53[8]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779__i8.GSR = "DISABLED";
    LUT4 i13250_2_lut_3_lut (.A(n18662), .B(n18586), .C(n153[3]), .Z(n199[3])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13250_2_lut_3_lut.init = 16'h7070;
    FD1P3IX SLO__i36 (.D(SLO[34]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i36.GSR = "DISABLED";
    FD1S3AX prev_MA_Temp_487 (.D(MA_Temp), .CK(clk), .Q(prev_MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam prev_MA_Temp_487.GSR = "DISABLED";
    FD1S3AX prev_MA_489 (.D(n30098), .CK(clk), .Q(prev_MA)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam prev_MA_489.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1779__i7 (.D(n53[7]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779__i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i0 (.D(\spi_data_out_r_39__N_4419[0] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i0.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1779__i6 (.D(n53[6]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779__i6.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1779__i5 (.D(n53[5]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779__i5.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1779__i4 (.D(n53[4]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779__i4.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1779__i3 (.D(n53[3]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779__i3.GSR = "DISABLED";
    LUT4 i13251_2_lut_3_lut (.A(n18662), .B(n18586), .C(n153[2]), .Z(n199[2])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13251_2_lut_3_lut.init = 16'h7070;
    FD1P3AX Cnt_NSL_1779__i2 (.D(n53[2]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779__i2.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1779__i1 (.D(n53[1]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779__i1.GSR = "DISABLED";
    LUT4 i24139_2_lut_3_lut_4_lut (.A(mode[2]), .B(n30103), .C(n30098), 
         .D(prev_MA), .Z(n12287)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i24139_2_lut_3_lut_4_lut.init = 16'h0020;
    FD1P3IX SLO__i15 (.D(SLO[13]), .SP(clk_enable_1120), .CD(GND_net), 
            .CK(clk), .Q(SLO[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i15.GSR = "DISABLED";
    LUT4 i13252_2_lut_3_lut (.A(n18662), .B(n18586), .C(n153[1]), .Z(n199[1])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13252_2_lut_3_lut.init = 16'h7070;
    LUT4 i24120_4_lut_4_lut (.A(mode[2]), .B(n30103), .C(n26373), .D(n30038), 
         .Z(clk_enable_1120)) /* synthesis lut_function=(!(A (B+(D))+!A ((D)+!C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i24120_4_lut_4_lut.init = 16'h0072;
    LUT4 i14110_3_lut_4_lut (.A(n30108), .B(n30107), .C(resetn_c), .D(n18586), 
         .Z(clk_1MHz_enable_70)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i14110_3_lut_4_lut.init = 16'h70f0;
    LUT4 n18662_bdd_3_lut (.A(n30034), .B(MA_Temp), .C(Cnt[5]), .Z(n29611)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam n18662_bdd_3_lut.init = 16'hc9c9;
    FD1P3IX mode__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_759), .CD(n30185), 
            .CK(clk), .Q(mode[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i0.GSR = "DISABLED";
    FD1P3IX SLO__i16 (.D(SLO[14]), .SP(clk_enable_1120), .CD(GND_net), 
            .CK(clk), .Q(SLO[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i16.GSR = "DISABLED";
    FD1P3IX SLO__i17 (.D(SLO[15]), .SP(clk_enable_1120), .CD(GND_net), 
            .CK(clk), .Q(SLO[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i17.GSR = "DISABLED";
    FD1P3IX SLO__i18 (.D(SLO[16]), .SP(clk_enable_1120), .CD(GND_net), 
            .CK(clk), .Q(SLO[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i18.GSR = "DISABLED";
    FD1P3IX SLO__i19 (.D(SLO[17]), .SP(clk_enable_1120), .CD(GND_net), 
            .CK(clk), .Q(SLO[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i19.GSR = "DISABLED";
    FD1P3IX SLO__i20 (.D(SLO[18]), .SP(clk_enable_1120), .CD(GND_net), 
            .CK(clk), .Q(SLO[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i20.GSR = "DISABLED";
    FD1P3AX SLO_buf__i1 (.D(SLO[0]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i1.GSR = "DISABLED";
    LUT4 n18662_bdd_4_lut (.A(n18662), .B(n30034), .C(MA_Temp), .D(Cnt[5]), 
         .Z(n29610)) /* synthesis lut_function=(!(A+!(B (C)+!B !(C (D)+!C !(D))))) */ ;
    defparam n18662_bdd_4_lut.init = 16'h4150;
    FD1S3IX spi_data_out_r_i39 (.D(\SLO_buf[13] ), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i39.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i38 (.D(\SLO_buf[12] ), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i38.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i37 (.D(\SLO_buf[11] ), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i37.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i36 (.D(\SLO_buf[10] ), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i36.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i35 (.D(\spi_data_out_r_39__N_4419[35] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i35.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i34 (.D(\spi_data_out_r_39__N_4419[34] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i34.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i33 (.D(\spi_data_out_r_39__N_4419[33] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i33.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_4419[32] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i31 (.D(SLO_buf[45]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i30 (.D(SLO_buf[44]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i29 (.D(SLO_buf[43]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i28 (.D(SLO_buf[42]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i27 (.D(SLO_buf[41]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i26 (.D(SLO_buf[40]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i25 (.D(SLO_buf[39]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i24 (.D(SLO_buf[38]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i23 (.D(SLO_buf[37]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i22 (.D(SLO_buf[36]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i21 (.D(SLO_buf[35]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i20 (.D(SLO_buf[34]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i19 (.D(SLO_buf[33]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i18 (.D(SLO_buf[32]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i17 (.D(SLO_buf[31]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i16 (.D(SLO_buf[30]), .CK(clk), .CD(n29992), 
            .Q(spi_data_out_r_39__N_4168[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_4419[15] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_4419[14] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_4419[13] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_4419[12] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_4419[11] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_4419[10] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_4419[9] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_4419[8] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_4419[7] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_4419[6] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_4419[5] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_4419[4] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_4419[3] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_4419[2] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_4419[1] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4168[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(\quad_homing[0] ), .B(pin_io_c_14), .Z(n25877)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(74[8:17])
    defparam i1_2_lut.init = 16'h8888;
    FD1S3IX i168_494 (.D(spi_data_out_r_39__N_4505), .CK(clk), .CD(n30185), 
            .Q(spi_data_out_r_39__N_4208)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam i168_494.GSR = "DISABLED";
    FD1P3IX digital_output_r_492 (.D(n28555), .SP(clk_enable_256), .CD(n30185), 
            .CK(clk), .Q(digital_output_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam digital_output_r_492.GSR = "DISABLED";
    FD1P3IX Cnt__i7 (.D(n199[7]), .SP(clk_1MHz_enable_41), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i7.GSR = "DISABLED";
    FD1P3IX Cnt__i6 (.D(n199[6]), .SP(clk_1MHz_enable_41), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i6.GSR = "DISABLED";
    FD1P3IX Cnt__i5 (.D(n199[5]), .SP(clk_1MHz_enable_41), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i5.GSR = "DISABLED";
    FD1P3IX Cnt__i4 (.D(n199[4]), .SP(clk_1MHz_enable_41), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i4.GSR = "DISABLED";
    FD1P3IX Cnt__i3 (.D(n199[3]), .SP(clk_1MHz_enable_41), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i3.GSR = "DISABLED";
    FD1P3IX Cnt__i2 (.D(n199[2]), .SP(clk_1MHz_enable_41), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i1 (.D(n199[1]), .SP(clk_1MHz_enable_41), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i1.GSR = "DISABLED";
    LUT4 i2972_2_lut_4_lut (.A(mode[2]), .B(mode[0]), .C(mode[1]), .D(pin_io_c_18), 
         .Z(\quad_a[1] )) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(107[27:54])
    defparam i2972_2_lut_4_lut.init = 16'h0400;
    LUT4 i2973_2_lut_4_lut (.A(mode[2]), .B(mode[0]), .C(mode[1]), .D(pin_io_out_19), 
         .Z(\quad_b[1] )) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(107[27:54])
    defparam i2973_2_lut_4_lut.init = 16'h0400;
    FD1P3IX MA_Temp_483 (.D(MA_Temp_N_4487), .SP(clk_1MHz_enable_42), .CD(n30185), 
            .CK(clk_1MHz), .Q(MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam MA_Temp_483.GSR = "DISABLED";
    FD1P3IX SLO__i2 (.D(SLO[0]), .SP(clk_enable_1120), .CD(GND_net), .CK(clk), 
            .Q(SLO[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i2.GSR = "DISABLED";
    FD1P3IX SLO__i3 (.D(SLO[1]), .SP(clk_enable_1120), .CD(GND_net), .CK(clk), 
            .Q(SLO[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i3.GSR = "DISABLED";
    FD1P3IX SLO__i4 (.D(SLO[2]), .SP(clk_enable_1120), .CD(GND_net), .CK(clk), 
            .Q(SLO[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i4.GSR = "DISABLED";
    FD1P3IX SLO__i5 (.D(SLO[3]), .SP(clk_enable_1120), .CD(GND_net), .CK(clk), 
            .Q(SLO[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i5.GSR = "DISABLED";
    FD1P3IX SLO__i21 (.D(SLO[19]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i21.GSR = "DISABLED";
    FD1P3IX SLO__i22 (.D(SLO[20]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i22.GSR = "DISABLED";
    FD1P3IX SLO__i37 (.D(SLO[35]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i37.GSR = "DISABLED";
    FD1P3IX SLO__i23 (.D(SLO[21]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i23.GSR = "DISABLED";
    FD1P3IX SLO__i24 (.D(SLO[22]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i24.GSR = "DISABLED";
    FD1P3IX SLO__i25 (.D(SLO[23]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i25.GSR = "DISABLED";
    FD1P3IX SLO__i38 (.D(SLO[36]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i38.GSR = "DISABLED";
    FD1P3IX SLO__i39 (.D(SLO[37]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i39.GSR = "DISABLED";
    FD1P3IX SLO__i40 (.D(SLO[38]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i40.GSR = "DISABLED";
    FD1P3IX SLO__i26 (.D(SLO[24]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i26.GSR = "DISABLED";
    FD1P3IX SLO__i27 (.D(SLO[25]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i27.GSR = "DISABLED";
    FD1P3IX SLO__i41 (.D(SLO[39]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i41.GSR = "DISABLED";
    FD1P3IX SLO__i42 (.D(SLO[40]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i42.GSR = "DISABLED";
    LUT4 i57_3_lut_4_lut (.A(mode[2]), .B(n30103), .C(uart_slot_en[0]), 
         .D(n30095), .Z(n28)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam i57_3_lut_4_lut.init = 16'hfe0e;
    FD1P3IX SLO__i28 (.D(SLO[26]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i28.GSR = "DISABLED";
    FD1P3IX mode__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_759), .CD(n30185), 
            .CK(clk), .Q(mode[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i1.GSR = "DISABLED";
    FD1P3IX mode__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_759), .CD(n30185), 
            .CK(clk), .Q(mode[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i2.GSR = "DISABLED";
    FD1P3IX SLO__i29 (.D(SLO[27]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i29.GSR = "DISABLED";
    FD1P3IX SLO__i30 (.D(SLO[28]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i30.GSR = "DISABLED";
    FD1P3AX SLO_buf__i2 (.D(SLO[1]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i2.GSR = "DISABLED";
    FD1P3IX SLO__i43 (.D(SLO[41]), .SP(clk_enable_1120), .CD(n12287), 
            .CK(clk), .Q(SLO[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i43.GSR = "DISABLED";
    FD1P3AX SLO_buf__i3 (.D(SLO[2]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i3.GSR = "DISABLED";
    FD1P3AX SLO_buf__i4 (.D(SLO[3]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i4.GSR = "DISABLED";
    FD1P3AX SLO_buf__i5 (.D(SLO[4]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i5.GSR = "DISABLED";
    FD1P3AX SLO_buf__i6 (.D(SLO[5]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i6.GSR = "DISABLED";
    FD1P3AX SLO_buf__i7 (.D(SLO[6]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i7.GSR = "DISABLED";
    FD1P3AX SLO_buf__i8 (.D(SLO[7]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i8.GSR = "DISABLED";
    FD1P3AX SLO_buf__i9 (.D(SLO[8]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i9.GSR = "DISABLED";
    FD1P3AX SLO_buf__i10 (.D(SLO[9]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i10.GSR = "DISABLED";
    FD1P3AX SLO_buf__i11 (.D(SLO[10]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i11.GSR = "DISABLED";
    FD1P3AX SLO_buf__i12 (.D(SLO[11]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i12.GSR = "DISABLED";
    FD1P3AX SLO_buf__i13 (.D(SLO[12]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i13.GSR = "DISABLED";
    FD1P3AX SLO_buf__i14 (.D(SLO[13]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i14.GSR = "DISABLED";
    FD1P3AX SLO_buf__i15 (.D(SLO[14]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i15.GSR = "DISABLED";
    FD1P3AX SLO_buf__i16 (.D(SLO[15]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i16.GSR = "DISABLED";
    FD1P3AX SLO_buf__i17 (.D(SLO[16]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i17.GSR = "DISABLED";
    FD1P3AX SLO_buf__i18 (.D(SLO[17]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i18.GSR = "DISABLED";
    FD1P3AX SLO_buf__i19 (.D(SLO[18]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i19.GSR = "DISABLED";
    FD1P3AX SLO_buf__i20 (.D(SLO[19]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i20.GSR = "DISABLED";
    FD1P3AX SLO_buf__i21 (.D(SLO[20]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i21.GSR = "DISABLED";
    FD1P3AX SLO_buf__i22 (.D(SLO[21]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i22.GSR = "DISABLED";
    FD1P3AX SLO_buf__i23 (.D(SLO[22]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i23.GSR = "DISABLED";
    FD1P3AX SLO_buf__i24 (.D(SLO[23]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i24.GSR = "DISABLED";
    FD1P3AX SLO_buf__i25 (.D(SLO[24]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i25.GSR = "DISABLED";
    FD1P3AX SLO_buf__i26 (.D(SLO[25]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i26.GSR = "DISABLED";
    FD1P3AX SLO_buf__i27 (.D(SLO[26]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i27.GSR = "DISABLED";
    FD1P3AX SLO_buf__i28 (.D(SLO[27]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i28.GSR = "DISABLED";
    FD1P3AX SLO_buf__i29 (.D(SLO[28]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i29.GSR = "DISABLED";
    FD1P3AX SLO_buf__i30 (.D(SLO[29]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(\SLO_buf[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i30.GSR = "DISABLED";
    FD1P3AX SLO_buf__i31 (.D(SLO[30]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i31.GSR = "DISABLED";
    FD1P3AX SLO_buf__i32 (.D(SLO[31]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i32.GSR = "DISABLED";
    FD1P3AX SLO_buf__i33 (.D(SLO[32]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i33.GSR = "DISABLED";
    FD1P3AX SLO_buf__i34 (.D(SLO[33]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i34.GSR = "DISABLED";
    FD1P3AX SLO_buf__i35 (.D(SLO[34]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i35.GSR = "DISABLED";
    FD1P3AX SLO_buf__i36 (.D(SLO[35]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i36.GSR = "DISABLED";
    FD1P3AX SLO_buf__i37 (.D(SLO[36]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i37.GSR = "DISABLED";
    FD1P3AX SLO_buf__i38 (.D(SLO[37]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i38.GSR = "DISABLED";
    FD1P3AX SLO_buf__i39 (.D(SLO[38]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i39.GSR = "DISABLED";
    FD1P3AX SLO_buf__i40 (.D(SLO[39]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i40.GSR = "DISABLED";
    FD1P3AX SLO_buf__i41 (.D(SLO[40]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i41.GSR = "DISABLED";
    FD1P3AX SLO_buf__i42 (.D(SLO[41]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i42.GSR = "DISABLED";
    FD1P3AX SLO_buf__i43 (.D(SLO[42]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i43.GSR = "DISABLED";
    FD1P3AX SLO_buf__i44 (.D(SLO[43]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i44.GSR = "DISABLED";
    FD1P3AX SLO_buf__i45 (.D(SLO[44]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i45.GSR = "DISABLED";
    FD1P3AX SLO_buf__i46 (.D(SLO[45]), .SP(SLO_buf_51__N_4358), .CK(clk), 
            .Q(SLO_buf[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i46.GSR = "DISABLED";
    FD1P3IX SLO__i6 (.D(SLO[4]), .SP(clk_enable_1120), .CD(GND_net), .CK(clk), 
            .Q(SLO[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i6.GSR = "DISABLED";
    LUT4 i23959_4_lut (.A(NSL), .B(n30042), .C(n18586), .D(n10368), 
         .Z(NSL_N_4500)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C+(D))))) */ ;
    defparam i23959_4_lut.init = 16'h3b37;
    FD1P3IX SLO__i7 (.D(SLO[5]), .SP(clk_enable_1120), .CD(GND_net), .CK(clk), 
            .Q(SLO[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i7.GSR = "DISABLED";
    LUT4 SLO_buf_51__I_118_2_lut (.A(prev_MA_Temp), .B(MA_Temp), .Z(SLO_buf_51__N_4358)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[5:38])
    defparam SLO_buf_51__I_118_2_lut.init = 16'h2222;
    FD1P3IX SLO__i8 (.D(SLO[6]), .SP(clk_enable_1120), .CD(GND_net), .CK(clk), 
            .Q(SLO[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i8.GSR = "DISABLED";
    LUT4 i23963_2_lut_rep_698 (.A(MA_Temp), .B(clk_1MHz), .Z(n30098)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i23963_2_lut_rep_698.init = 16'h7777;
    PFUMX i24281 (.BLUT(n29611), .ALUT(n29610), .C0(n18586), .Z(MA_Temp_N_4487));
    LUT4 i1_2_lut_rep_638_3_lut (.A(MA_Temp), .B(clk_1MHz), .C(prev_MA), 
         .Z(n30038)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i1_2_lut_rep_638_3_lut.init = 16'hf8f8;
    LUT4 digital_output_r_I_0_547_3_lut (.A(digital_output_r), .B(UC_TXD0_c), 
         .C(OW_ID_N_4462), .Z(OW_ID_N_4461)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[16] 91[59])
    defparam digital_output_r_I_0_547_3_lut.init = 16'hcaca;
    LUT4 i24066_4_lut (.A(OW_ID_N_4462), .B(mode[1]), .C(mode[0]), .D(mode[2]), 
         .Z(OW_ID_N_4467)) /* synthesis lut_function=(!(A+!((C+(D))+!B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[8:13])
    defparam i24066_4_lut.init = 16'h5551;
    LUT4 i5_3_lut (.A(mode[1]), .B(n10_adj_6707), .C(uart_slot_en[0]), 
         .Z(OW_ID_N_4462)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i5_3_lut.init = 16'h0404;
    LUT4 i4_4_lut (.A(mode[0]), .B(n30050), .C(mode[2]), .D(uart_slot_en[1]), 
         .Z(n10_adj_6707)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i4_4_lut.init = 16'h0008;
    CCU2D add_564_9 (.A0(Cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21927), 
          .S0(n153[7]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_9.INIT0 = 16'h5aaa;
    defparam add_564_9.INIT1 = 16'h0000;
    defparam add_564_9.INJECT1_0 = "NO";
    defparam add_564_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_703 (.A(mode[0]), .B(mode[1]), .Z(n30103)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_rep_703.init = 16'heeee;
    LUT4 i1_2_lut_rep_641_3_lut (.A(mode[0]), .B(mode[1]), .C(mode[2]), 
         .Z(n30041)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_rep_641_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_4_lut (.A(mode[0]), .B(mode[1]), .C(Cnt[5]), .D(mode[2]), 
         .Z(n26297)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfeff;
    LUT4 i1_2_lut_rep_675_3_lut (.A(mode[0]), .B(mode[1]), .C(mode[2]), 
         .Z(n30075)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_rep_675_3_lut.init = 16'hfefe;
    LUT4 i2970_2_lut_3_lut_4_lut (.A(mode[0]), .B(mode[1]), .C(pin_io_c_13), 
         .D(mode[2]), .Z(\pin_intrpt[4] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2970_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 RESET_N_4460_bdd_2_lut_3_lut_4_lut (.A(mode[0]), .B(mode[1]), .C(pin_io_out_15), 
         .D(mode[2]), .Z(n29944)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam RESET_N_4460_bdd_2_lut_3_lut_4_lut.init = 16'hf0e0;
    CCU2D add_564_7 (.A0(Cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21926), 
          .COUT(n21927), .S0(n153[5]), .S1(n153[6]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_7.INIT0 = 16'h5aaa;
    defparam add_564_7.INIT1 = 16'h5aaa;
    defparam add_564_7.INJECT1_0 = "NO";
    defparam add_564_7.INJECT1_1 = "NO";
    LUT4 i2969_2_lut_3_lut_4_lut (.A(mode[0]), .B(mode[1]), .C(pin_io_c_12), 
         .D(mode[2]), .Z(\pin_intrpt[3] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2969_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2971_2_lut_3_lut_4_lut (.A(mode[0]), .B(mode[1]), .C(pin_io_c_14), 
         .D(mode[2]), .Z(\pin_intrpt[5] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2971_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2963_1_lut_2_lut_3_lut (.A(mode[0]), .B(mode[1]), .C(mode[2]), 
         .Z(n7277)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2963_1_lut_2_lut_3_lut.init = 16'h0101;
    LUT4 i23926_2_lut_3_lut_4_lut (.A(n30042), .B(resetn_c), .C(n18586), 
         .D(n18662), .Z(clk_1MHz_enable_42)) /* synthesis lut_function=(!(A (C (D))+!A (B+(C (D))))) */ ;
    defparam i23926_2_lut_3_lut_4_lut.init = 16'h0bbb;
    LUT4 i2442_2_lut_rep_704 (.A(mode[0]), .B(mode[1]), .Z(n30104)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2442_2_lut_rep_704.init = 16'h8888;
    LUT4 i24069_2_lut_3_lut (.A(mode[0]), .B(mode[1]), .C(mode[2]), .Z(ENC_O_N_4469)) /* synthesis lut_function=(!(A (B+(C))+!A (C))) */ ;
    defparam i24069_2_lut_3_lut.init = 16'h0707;
    LUT4 i1_2_lut_rep_705 (.A(Cnt[7]), .B(Cnt[6]), .Z(n30105)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_705.init = 16'heeee;
    LUT4 i1_3_lut_4_lut (.A(Cnt[7]), .B(Cnt[6]), .C(Cnt[0]), .D(n30106), 
         .Z(n11629)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hfffe;
    LUT4 i12925_2_lut_3_lut (.A(n18662), .B(n18586), .C(n153[0]), .Z(n199[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i12925_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_706 (.A(Cnt[2]), .B(Cnt[3]), .Z(n30106)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(109[8:17])
    defparam i1_2_lut_rep_706.init = 16'heeee;
    LUT4 i13246_2_lut_3_lut (.A(n18662), .B(n18586), .C(n153[7]), .Z(n199[7])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13246_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_3_lut_4_lut_adj_590 (.A(Cnt[2]), .B(Cnt[3]), .C(Cnt[1]), .D(Cnt[0]), 
         .Z(n18478)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(109[8:17])
    defparam i1_3_lut_4_lut_adj_590.init = 16'hfeee;
    LUT4 i1_3_lut_rep_707 (.A(Cnt_NSL[9]), .B(Cnt_NSL[8]), .C(Cnt_NSL[7]), 
         .Z(n30107)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_rep_707.init = 16'hfefe;
    LUT4 i1_2_lut_rep_642_4_lut (.A(Cnt_NSL[9]), .B(Cnt_NSL[8]), .C(Cnt_NSL[7]), 
         .D(n30108), .Z(n30042)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_rep_642_4_lut.init = 16'hfe00;
    CCU2D add_564_5 (.A0(Cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21925), 
          .COUT(n21926), .S0(n153[3]), .S1(n153[4]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_5.INIT0 = 16'h5aaa;
    defparam add_564_5.INIT1 = 16'h5aaa;
    defparam add_564_5.INJECT1_0 = "NO";
    defparam add_564_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_708 (.A(Cnt_NSL[11]), .B(Cnt_NSL[10]), .Z(n30108)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i1_2_lut_rep_708.init = 16'h8888;
    LUT4 i24028_2_lut_rep_614_3_lut_4_lut (.A(Cnt_NSL[11]), .B(Cnt_NSL[10]), 
         .C(resetn_c), .D(n30107), .Z(clk_1MHz_enable_41)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i24028_2_lut_rep_614_3_lut_4_lut.init = 16'h8f0f;
    CCU2D add_564_3 (.A0(Cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21924), 
          .COUT(n21925), .S0(n153[1]), .S1(n153[2]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_3.INIT0 = 16'h5aaa;
    defparam add_564_3.INIT1 = 16'h5aaa;
    defparam add_564_3.INJECT1_0 = "NO";
    defparam add_564_3.INJECT1_1 = "NO";
    LUT4 i13247_2_lut_3_lut (.A(n18662), .B(n18586), .C(n153[6]), .Z(n199[6])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13247_2_lut_3_lut.init = 16'h7070;
    LUT4 i13248_2_lut_3_lut (.A(n18662), .B(n18586), .C(n153[5]), .Z(n199[5])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13248_2_lut_3_lut.init = 16'h7070;
    CCU2D add_564_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n21924), 
          .S1(n153[0]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_1.INIT0 = 16'hF000;
    defparam add_564_1.INIT1 = 16'h5555;
    defparam add_564_1.INJECT1_0 = "NO";
    defparam add_564_1.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1779_add_4_13 (.A0(Cnt_NSL[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21923), .S0(n53[11]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779_add_4_13.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1779_add_4_13.INIT1 = 16'h0000;
    defparam Cnt_NSL_1779_add_4_13.INJECT1_0 = "NO";
    defparam Cnt_NSL_1779_add_4_13.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1779_add_4_11 (.A0(Cnt_NSL[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Cnt_NSL[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21922), .COUT(n21923), .S0(n53[9]), .S1(n53[10]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779_add_4_11.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1779_add_4_11.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1779_add_4_11.INJECT1_0 = "NO";
    defparam Cnt_NSL_1779_add_4_11.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1779_add_4_9 (.A0(Cnt_NSL[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Cnt_NSL[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n21921), .COUT(n21922), .S0(n53[7]), .S1(n53[8]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779_add_4_9.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1779_add_4_9.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1779_add_4_9.INJECT1_0 = "NO";
    defparam Cnt_NSL_1779_add_4_9.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1779_add_4_7 (.A0(n93[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21920), .COUT(n21921), .S0(n53[5]), .S1(n53[6]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779_add_4_7.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1779_add_4_7.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1779_add_4_7.INJECT1_0 = "NO";
    defparam Cnt_NSL_1779_add_4_7.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1779_add_4_5 (.A0(n93[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21919), .COUT(n21920), .S0(n53[3]), .S1(n53[4]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779_add_4_5.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1779_add_4_5.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1779_add_4_5.INJECT1_0 = "NO";
    defparam Cnt_NSL_1779_add_4_5.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1779_add_4_3 (.A0(n93[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n21918), .COUT(n21919), .S0(n53[1]), .S1(n53[2]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779_add_4_3.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1779_add_4_3.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1779_add_4_3.INJECT1_0 = "NO";
    defparam Cnt_NSL_1779_add_4_3.INJECT1_1 = "NO";
    FD1P3AX NSL_484 (.D(NSL_N_4500), .SP(clk_1MHz_enable_70), .CK(clk_1MHz), 
            .Q(NSL)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam NSL_484.GSR = "DISABLED";
    FD1P3IX SLO__i9 (.D(SLO[7]), .SP(clk_enable_1120), .CD(GND_net), .CK(clk), 
            .Q(SLO[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i9.GSR = "DISABLED";
    FD1P3IX SLO__i10 (.D(SLO[8]), .SP(clk_enable_1120), .CD(GND_net), 
            .CK(clk), .Q(SLO[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i10.GSR = "DISABLED";
    CCU2D Cnt_NSL_1779_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n30107), .B1(n30108), .C1(n93[0]), .D1(GND_net), 
          .COUT(n21918), .S1(n53[0]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1779_add_4_1.INIT0 = 16'hF000;
    defparam Cnt_NSL_1779_add_4_1.INIT1 = 16'h8787;
    defparam Cnt_NSL_1779_add_4_1.INJECT1_0 = "NO";
    defparam Cnt_NSL_1779_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_718 (.A(UC_TXD0_c), .B(uart_slot_en[3]), .Z(n30118)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_rep_718.init = 16'h4444;
    FD1P3IX SLO__i11 (.D(SLO[9]), .SP(clk_enable_1120), .CD(GND_net), 
            .CK(clk), .Q(SLO[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i11.GSR = "DISABLED";
    LUT4 i2_3_lut_rep_649_4_lut (.A(UC_TXD0_c), .B(uart_slot_en[3]), .C(uart_slot_en[2]), 
         .D(uart_slot_en[1]), .Z(n30049)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i2_3_lut_rep_649_4_lut.init = 16'h0040;
    LUT4 i2_2_lut_rep_650_3_lut (.A(UC_TXD0_c), .B(uart_slot_en[3]), .C(uart_slot_en[2]), 
         .Z(n30050)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i2_2_lut_rep_650_3_lut.init = 16'h0404;
    LUT4 i3_2_lut_3_lut_4_lut (.A(UC_TXD0_c), .B(uart_slot_en[3]), .C(\mode[2] ), 
         .D(uart_slot_en[2]), .Z(n9)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i3_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i1_4_lut (.A(n30105), .B(n25214), .C(n30104), .D(mode[2]), 
         .Z(n18662)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i1_4_lut.init = 16'hffef;
    LUT4 i1_3_lut (.A(Cnt[5]), .B(n18478), .C(Cnt[4]), .Z(n25214)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_adj_591 (.A(n30105), .B(n18478), .C(n26297), .D(Cnt[4]), 
         .Z(n18586)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_591.init = 16'hfefa;
    LUT4 i1_3_lut_adj_592 (.A(mode[1]), .B(mode[0]), .C(n24765), .Z(n26373)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_592.init = 16'h8080;
    LUT4 i3_4_lut (.A(Cnt[5]), .B(Cnt[1]), .C(n11629), .D(Cnt[4]), .Z(n24765)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(133[16:19])
    defparam i3_4_lut.init = 16'hfffe;
    
endmodule
//
// Verilog Description of module \quad_decoder(DEV_ID=2) 
//

module \quad_decoder(DEV_ID=2)  (quad_homing, clk, clk_enable_488, n30185, 
            \spi_data_r[0] , quad_count, \quad_b[2] , \spi_data_out_r_39__N_1404[0] , 
            \spi_data_out_r_39__N_1553[0] , quad_buffer, \pin_intrpt[8] , 
            clk_enable_211, \quad_a[2] , \spi_data_r[31] , \spi_data_r[30] , 
            \spi_data_r[29] , \spi_data_r[28] , \spi_data_r[27] , \spi_data_r[26] , 
            \spi_data_r[25] , \spi_data_r[24] , \spi_data_r[23] , \spi_data_r[22] , 
            \spi_data_r[21] , \spi_data_r[20] , \spi_data_r[19] , \spi_data_r[18] , 
            \spi_data_r[17] , \spi_data_r[16] , \spi_data_r[15] , \spi_data_r[14] , 
            \spi_data_r[13] , \spi_data_r[12] , \spi_data_r[11] , \spi_data_r[10] , 
            \spi_data_r[9] , \spi_data_r[8] , \spi_data_r[7] , \spi_data_r[6] , 
            \spi_data_r[5] , \spi_data_r[4] , \spi_data_r[3] , \spi_data_r[2] , 
            \spi_data_r[1] , spi_data_out_r_39__N_1444, spi_data_out_r_39__N_1633, 
            n29993, \spi_data_out_r_39__N_1404[31] , \spi_data_out_r_39__N_1553[31] , 
            \spi_data_out_r_39__N_1404[30] , \spi_data_out_r_39__N_1553[30] , 
            \spi_data_out_r_39__N_1404[29] , \spi_data_out_r_39__N_1553[29] , 
            \spi_data_out_r_39__N_1404[28] , \spi_data_out_r_39__N_1553[28] , 
            \spi_data_out_r_39__N_1404[27] , \spi_data_out_r_39__N_1553[27] , 
            \spi_data_out_r_39__N_1404[26] , \spi_data_out_r_39__N_1553[26] , 
            \spi_data_out_r_39__N_1404[25] , \spi_data_out_r_39__N_1553[25] , 
            \spi_data_out_r_39__N_1404[24] , \spi_data_out_r_39__N_1553[24] , 
            \spi_data_out_r_39__N_1404[23] , \spi_data_out_r_39__N_1553[23] , 
            \spi_data_out_r_39__N_1404[22] , \spi_data_out_r_39__N_1553[22] , 
            \spi_data_out_r_39__N_1404[21] , \spi_data_out_r_39__N_1553[21] , 
            \spi_data_out_r_39__N_1404[20] , \spi_data_out_r_39__N_1553[20] , 
            \spi_data_out_r_39__N_1404[19] , \spi_data_out_r_39__N_1553[19] , 
            \spi_data_out_r_39__N_1404[18] , \spi_data_out_r_39__N_1553[18] , 
            \spi_data_out_r_39__N_1404[17] , \spi_data_out_r_39__N_1553[17] , 
            \spi_data_out_r_39__N_1404[16] , \spi_data_out_r_39__N_1553[16] , 
            \spi_data_out_r_39__N_1404[15] , \spi_data_out_r_39__N_1553[15] , 
            \spi_data_out_r_39__N_1404[14] , \spi_data_out_r_39__N_1553[14] , 
            \spi_data_out_r_39__N_1404[13] , \spi_data_out_r_39__N_1553[13] , 
            \spi_data_out_r_39__N_1404[12] , \spi_data_out_r_39__N_1553[12] , 
            \spi_data_out_r_39__N_1404[11] , \spi_data_out_r_39__N_1553[11] , 
            \spi_data_out_r_39__N_1404[10] , \spi_data_out_r_39__N_1553[10] , 
            \spi_data_out_r_39__N_1404[9] , \spi_data_out_r_39__N_1553[9] , 
            \spi_data_out_r_39__N_1404[8] , \spi_data_out_r_39__N_1553[8] , 
            \spi_data_out_r_39__N_1404[7] , \spi_data_out_r_39__N_1553[7] , 
            \spi_data_out_r_39__N_1404[6] , \spi_data_out_r_39__N_1553[6] , 
            \spi_data_out_r_39__N_1404[5] , \spi_data_out_r_39__N_1553[5] , 
            \spi_data_out_r_39__N_1404[4] , \spi_data_out_r_39__N_1553[4] , 
            \spi_data_out_r_39__N_1404[3] , \spi_data_out_r_39__N_1553[3] , 
            \spi_data_out_r_39__N_1404[2] , \spi_data_out_r_39__N_1553[2] , 
            \spi_data_out_r_39__N_1404[1] , \spi_data_out_r_39__N_1553[1] , 
            resetn_c, n1, GND_net) /* synthesis syn_module_defined=1 */ ;
    output [1:0]quad_homing;
    input clk;
    input clk_enable_488;
    input n30185;
    input \spi_data_r[0] ;
    output [31:0]quad_count;
    input \quad_b[2] ;
    output \spi_data_out_r_39__N_1404[0] ;
    input \spi_data_out_r_39__N_1553[0] ;
    output [31:0]quad_buffer;
    input \pin_intrpt[8] ;
    input clk_enable_211;
    input \quad_a[2] ;
    input \spi_data_r[31] ;
    input \spi_data_r[30] ;
    input \spi_data_r[29] ;
    input \spi_data_r[28] ;
    input \spi_data_r[27] ;
    input \spi_data_r[26] ;
    input \spi_data_r[25] ;
    input \spi_data_r[24] ;
    input \spi_data_r[23] ;
    input \spi_data_r[22] ;
    input \spi_data_r[21] ;
    input \spi_data_r[20] ;
    input \spi_data_r[19] ;
    input \spi_data_r[18] ;
    input \spi_data_r[17] ;
    input \spi_data_r[16] ;
    input \spi_data_r[15] ;
    input \spi_data_r[14] ;
    input \spi_data_r[13] ;
    input \spi_data_r[12] ;
    input \spi_data_r[11] ;
    input \spi_data_r[10] ;
    input \spi_data_r[9] ;
    input \spi_data_r[8] ;
    input \spi_data_r[7] ;
    input \spi_data_r[6] ;
    input \spi_data_r[5] ;
    input \spi_data_r[4] ;
    input \spi_data_r[3] ;
    input \spi_data_r[2] ;
    input \spi_data_r[1] ;
    output spi_data_out_r_39__N_1444;
    input spi_data_out_r_39__N_1633;
    input n29993;
    output \spi_data_out_r_39__N_1404[31] ;
    input \spi_data_out_r_39__N_1553[31] ;
    output \spi_data_out_r_39__N_1404[30] ;
    input \spi_data_out_r_39__N_1553[30] ;
    output \spi_data_out_r_39__N_1404[29] ;
    input \spi_data_out_r_39__N_1553[29] ;
    output \spi_data_out_r_39__N_1404[28] ;
    input \spi_data_out_r_39__N_1553[28] ;
    output \spi_data_out_r_39__N_1404[27] ;
    input \spi_data_out_r_39__N_1553[27] ;
    output \spi_data_out_r_39__N_1404[26] ;
    input \spi_data_out_r_39__N_1553[26] ;
    output \spi_data_out_r_39__N_1404[25] ;
    input \spi_data_out_r_39__N_1553[25] ;
    output \spi_data_out_r_39__N_1404[24] ;
    input \spi_data_out_r_39__N_1553[24] ;
    output \spi_data_out_r_39__N_1404[23] ;
    input \spi_data_out_r_39__N_1553[23] ;
    output \spi_data_out_r_39__N_1404[22] ;
    input \spi_data_out_r_39__N_1553[22] ;
    output \spi_data_out_r_39__N_1404[21] ;
    input \spi_data_out_r_39__N_1553[21] ;
    output \spi_data_out_r_39__N_1404[20] ;
    input \spi_data_out_r_39__N_1553[20] ;
    output \spi_data_out_r_39__N_1404[19] ;
    input \spi_data_out_r_39__N_1553[19] ;
    output \spi_data_out_r_39__N_1404[18] ;
    input \spi_data_out_r_39__N_1553[18] ;
    output \spi_data_out_r_39__N_1404[17] ;
    input \spi_data_out_r_39__N_1553[17] ;
    output \spi_data_out_r_39__N_1404[16] ;
    input \spi_data_out_r_39__N_1553[16] ;
    output \spi_data_out_r_39__N_1404[15] ;
    input \spi_data_out_r_39__N_1553[15] ;
    output \spi_data_out_r_39__N_1404[14] ;
    input \spi_data_out_r_39__N_1553[14] ;
    output \spi_data_out_r_39__N_1404[13] ;
    input \spi_data_out_r_39__N_1553[13] ;
    output \spi_data_out_r_39__N_1404[12] ;
    input \spi_data_out_r_39__N_1553[12] ;
    output \spi_data_out_r_39__N_1404[11] ;
    input \spi_data_out_r_39__N_1553[11] ;
    output \spi_data_out_r_39__N_1404[10] ;
    input \spi_data_out_r_39__N_1553[10] ;
    output \spi_data_out_r_39__N_1404[9] ;
    input \spi_data_out_r_39__N_1553[9] ;
    output \spi_data_out_r_39__N_1404[8] ;
    input \spi_data_out_r_39__N_1553[8] ;
    output \spi_data_out_r_39__N_1404[7] ;
    input \spi_data_out_r_39__N_1553[7] ;
    output \spi_data_out_r_39__N_1404[6] ;
    input \spi_data_out_r_39__N_1553[6] ;
    output \spi_data_out_r_39__N_1404[5] ;
    input \spi_data_out_r_39__N_1553[5] ;
    output \spi_data_out_r_39__N_1404[4] ;
    input \spi_data_out_r_39__N_1553[4] ;
    output \spi_data_out_r_39__N_1404[3] ;
    input \spi_data_out_r_39__N_1553[3] ;
    output \spi_data_out_r_39__N_1404[2] ;
    input \spi_data_out_r_39__N_1553[2] ;
    output \spi_data_out_r_39__N_1404[1] ;
    input \spi_data_out_r_39__N_1553[1] ;
    input resetn_c;
    input n1;
    input GND_net;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire \pin_intrpt[8]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[8] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    
    wire clk_enable_485, n7981;
    wire [2:0]quad_b_delayed;   // c:/s_links/sources/quad_decoder.v(35[19:33])
    wire [31:0]quad_set;   // c:/s_links/sources/quad_decoder.v(39[31:39])
    wire [2:0]quad_a_delayed;   // c:/s_links/sources/quad_decoder.v(34[20:34])
    
    wire n22105, n6;
    wire [31:0]n4063;
    
    wire n22104, n22103, n22102, n22101, quad_set_valid, n22100, 
        n22099, n22098, n22097, n22096, n22095, n22094, n22093, 
        n8648, n8650, n8652, n8654, n8656, n8658, n8660, n8662, 
        n8664, n8666, n8668, n8670, n8672, n8674, n8676, n8678, 
        n8680, n8682, n8684, n8686, n8688, n8690, n8692, n8694, 
        n8696, n8698, n8700, n8702, n8704, n8706, n8708, n22092, 
        n22091, n5703, n22090, count_dir;
    
    FD1P3IX quad_homing__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_488), .CD(n30185), 
            .CK(clk), .Q(quad_homing[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(62[8] 69[4])
    defparam quad_homing__i0.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i0 (.D(n7981), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i0.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i0 (.D(\quad_b[2] ), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_1553[0] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX quad_buffer_i0 (.D(quad_count[0]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i0.GSR = "DISABLED";
    FD1P3IX quad_set__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i0.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i0 (.D(\quad_a[2] ), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i0.GSR = "DISABLED";
    FD1P3IX quad_set__i31 (.D(\spi_data_r[31] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i31.GSR = "DISABLED";
    FD1P3IX quad_set__i30 (.D(\spi_data_r[30] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i30.GSR = "DISABLED";
    FD1P3IX quad_set__i29 (.D(\spi_data_r[29] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i29.GSR = "DISABLED";
    FD1P3IX quad_set__i28 (.D(\spi_data_r[28] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i28.GSR = "DISABLED";
    FD1P3IX quad_set__i27 (.D(\spi_data_r[27] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i27.GSR = "DISABLED";
    FD1P3IX quad_set__i26 (.D(\spi_data_r[26] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i26.GSR = "DISABLED";
    FD1P3IX quad_set__i25 (.D(\spi_data_r[25] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i25.GSR = "DISABLED";
    FD1P3IX quad_set__i24 (.D(\spi_data_r[24] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i24.GSR = "DISABLED";
    FD1P3IX quad_set__i23 (.D(\spi_data_r[23] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i23.GSR = "DISABLED";
    FD1P3IX quad_set__i22 (.D(\spi_data_r[22] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i22.GSR = "DISABLED";
    FD1P3IX quad_set__i21 (.D(\spi_data_r[21] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i21.GSR = "DISABLED";
    FD1P3IX quad_set__i20 (.D(\spi_data_r[20] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i20.GSR = "DISABLED";
    FD1P3IX quad_set__i19 (.D(\spi_data_r[19] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i19.GSR = "DISABLED";
    FD1P3IX quad_set__i18 (.D(\spi_data_r[18] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i18.GSR = "DISABLED";
    FD1P3IX quad_set__i17 (.D(\spi_data_r[17] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i17.GSR = "DISABLED";
    FD1P3IX quad_set__i16 (.D(\spi_data_r[16] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i16.GSR = "DISABLED";
    FD1P3IX quad_set__i15 (.D(\spi_data_r[15] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i15.GSR = "DISABLED";
    FD1P3IX quad_set__i14 (.D(\spi_data_r[14] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i14.GSR = "DISABLED";
    FD1P3IX quad_set__i13 (.D(\spi_data_r[13] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i13.GSR = "DISABLED";
    FD1P3IX quad_set__i12 (.D(\spi_data_r[12] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i12.GSR = "DISABLED";
    FD1P3IX quad_set__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i11.GSR = "DISABLED";
    FD1P3IX quad_set__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i10.GSR = "DISABLED";
    FD1P3IX quad_set__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i9.GSR = "DISABLED";
    FD1P3IX quad_set__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i8.GSR = "DISABLED";
    FD1P3IX quad_set__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i7.GSR = "DISABLED";
    FD1P3IX quad_set__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i6.GSR = "DISABLED";
    FD1P3IX quad_set__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i5.GSR = "DISABLED";
    FD1P3IX quad_set__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i4.GSR = "DISABLED";
    FD1P3IX quad_set__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i3.GSR = "DISABLED";
    FD1P3IX quad_set__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i2.GSR = "DISABLED";
    FD1P3IX quad_set__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_211), .CD(n30185), 
            .CK(clk), .Q(quad_set[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i1.GSR = "DISABLED";
    CCU2D add_1365_33 (.A0(quad_count[30]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[31]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22105), .S0(n4063[30]), .S1(n4063[31]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_33.INIT0 = 16'h5569;
    defparam add_1365_33.INIT1 = 16'h5569;
    defparam add_1365_33.INJECT1_0 = "NO";
    defparam add_1365_33.INJECT1_1 = "NO";
    CCU2D add_1365_31 (.A0(quad_count[28]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[29]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22104), .COUT(n22105), .S0(n4063[28]), .S1(n4063[29]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_31.INIT0 = 16'h5569;
    defparam add_1365_31.INIT1 = 16'h5569;
    defparam add_1365_31.INJECT1_0 = "NO";
    defparam add_1365_31.INJECT1_1 = "NO";
    CCU2D add_1365_29 (.A0(quad_count[26]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[27]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22103), .COUT(n22104), .S0(n4063[26]), .S1(n4063[27]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_29.INIT0 = 16'h5569;
    defparam add_1365_29.INIT1 = 16'h5569;
    defparam add_1365_29.INJECT1_0 = "NO";
    defparam add_1365_29.INJECT1_1 = "NO";
    CCU2D add_1365_27 (.A0(quad_count[24]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[25]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22102), .COUT(n22103), .S0(n4063[24]), .S1(n4063[25]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_27.INIT0 = 16'h5569;
    defparam add_1365_27.INIT1 = 16'h5569;
    defparam add_1365_27.INJECT1_0 = "NO";
    defparam add_1365_27.INJECT1_1 = "NO";
    FD1S3IX i39_391 (.D(spi_data_out_r_39__N_1633), .CK(clk), .CD(n30185), 
            .Q(spi_data_out_r_39__N_1444)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam i39_391.GSR = "DISABLED";
    CCU2D add_1365_25 (.A0(quad_count[22]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[23]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22101), .COUT(n22102), .S0(n4063[22]), .S1(n4063[23]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_25.INIT0 = 16'h5569;
    defparam add_1365_25.INIT1 = 16'h5569;
    defparam add_1365_25.INJECT1_0 = "NO";
    defparam add_1365_25.INJECT1_1 = "NO";
    FD1S3IX quad_set_valid_388 (.D(n29993), .CK(clk), .CD(n30185), .Q(quad_set_valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set_valid_388.GSR = "DISABLED";
    CCU2D add_1365_23 (.A0(quad_count[20]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[21]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22100), .COUT(n22101), .S0(n4063[20]), .S1(n4063[21]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_23.INIT0 = 16'h5569;
    defparam add_1365_23.INIT1 = 16'h5569;
    defparam add_1365_23.INJECT1_0 = "NO";
    defparam add_1365_23.INJECT1_1 = "NO";
    CCU2D add_1365_21 (.A0(quad_count[18]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[19]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22099), .COUT(n22100), .S0(n4063[18]), .S1(n4063[19]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_21.INIT0 = 16'h5569;
    defparam add_1365_21.INIT1 = 16'h5569;
    defparam add_1365_21.INJECT1_0 = "NO";
    defparam add_1365_21.INJECT1_1 = "NO";
    CCU2D add_1365_19 (.A0(quad_count[16]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[17]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22098), .COUT(n22099), .S0(n4063[16]), .S1(n4063[17]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_19.INIT0 = 16'h5569;
    defparam add_1365_19.INIT1 = 16'h5569;
    defparam add_1365_19.INJECT1_0 = "NO";
    defparam add_1365_19.INJECT1_1 = "NO";
    CCU2D add_1365_17 (.A0(quad_count[14]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[15]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22097), .COUT(n22098), .S0(n4063[14]), .S1(n4063[15]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_17.INIT0 = 16'h5569;
    defparam add_1365_17.INIT1 = 16'h5569;
    defparam add_1365_17.INJECT1_0 = "NO";
    defparam add_1365_17.INJECT1_1 = "NO";
    CCU2D add_1365_15 (.A0(quad_count[12]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[13]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22096), .COUT(n22097), .S0(n4063[12]), .S1(n4063[13]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_15.INIT0 = 16'h5569;
    defparam add_1365_15.INIT1 = 16'h5569;
    defparam add_1365_15.INJECT1_0 = "NO";
    defparam add_1365_15.INJECT1_1 = "NO";
    CCU2D add_1365_13 (.A0(quad_count[10]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[11]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22095), .COUT(n22096), .S0(n4063[10]), .S1(n4063[11]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_13.INIT0 = 16'h5569;
    defparam add_1365_13.INIT1 = 16'h5569;
    defparam add_1365_13.INJECT1_0 = "NO";
    defparam add_1365_13.INJECT1_1 = "NO";
    CCU2D add_1365_11 (.A0(quad_count[8]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[9]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22094), .COUT(n22095), .S0(n4063[8]), .S1(n4063[9]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_11.INIT0 = 16'h5569;
    defparam add_1365_11.INIT1 = 16'h5569;
    defparam add_1365_11.INJECT1_0 = "NO";
    defparam add_1365_11.INJECT1_1 = "NO";
    CCU2D add_1365_9 (.A0(quad_count[6]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[7]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22093), .COUT(n22094), .S0(n4063[6]), .S1(n4063[7]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_9.INIT0 = 16'h5569;
    defparam add_1365_9.INIT1 = 16'h5569;
    defparam add_1365_9.INJECT1_0 = "NO";
    defparam add_1365_9.INJECT1_1 = "NO";
    FD1S3AX quad_buffer_i31 (.D(quad_count[31]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i31.GSR = "DISABLED";
    FD1S3AX quad_buffer_i30 (.D(quad_count[30]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i30.GSR = "DISABLED";
    FD1S3AX quad_buffer_i29 (.D(quad_count[29]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i29.GSR = "DISABLED";
    FD1S3AX quad_buffer_i28 (.D(quad_count[28]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i28.GSR = "DISABLED";
    FD1S3AX quad_buffer_i27 (.D(quad_count[27]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i27.GSR = "DISABLED";
    FD1S3AX quad_buffer_i26 (.D(quad_count[26]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i26.GSR = "DISABLED";
    FD1S3AX quad_buffer_i25 (.D(quad_count[25]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i25.GSR = "DISABLED";
    FD1S3AX quad_buffer_i24 (.D(quad_count[24]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i24.GSR = "DISABLED";
    FD1S3AX quad_buffer_i23 (.D(quad_count[23]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i23.GSR = "DISABLED";
    FD1S3AX quad_buffer_i22 (.D(quad_count[22]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i22.GSR = "DISABLED";
    FD1S3AX quad_buffer_i21 (.D(quad_count[21]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i21.GSR = "DISABLED";
    FD1S3AX quad_buffer_i20 (.D(quad_count[20]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i20.GSR = "DISABLED";
    FD1S3AX quad_buffer_i19 (.D(quad_count[19]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i19.GSR = "DISABLED";
    FD1S3AX quad_buffer_i18 (.D(quad_count[18]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i18.GSR = "DISABLED";
    FD1S3AX quad_buffer_i17 (.D(quad_count[17]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i17.GSR = "DISABLED";
    FD1S3AX quad_buffer_i16 (.D(quad_count[16]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i16.GSR = "DISABLED";
    FD1S3AX quad_buffer_i15 (.D(quad_count[15]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i15.GSR = "DISABLED";
    FD1S3AX quad_buffer_i14 (.D(quad_count[14]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i14.GSR = "DISABLED";
    FD1S3AX quad_buffer_i13 (.D(quad_count[13]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i13.GSR = "DISABLED";
    FD1S3AX quad_buffer_i12 (.D(quad_count[12]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i12.GSR = "DISABLED";
    FD1S3AX quad_buffer_i11 (.D(quad_count[11]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i11.GSR = "DISABLED";
    FD1S3AX quad_buffer_i10 (.D(quad_count[10]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i10.GSR = "DISABLED";
    FD1S3AX quad_buffer_i9 (.D(quad_count[9]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i9.GSR = "DISABLED";
    FD1S3AX quad_buffer_i8 (.D(quad_count[8]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i8.GSR = "DISABLED";
    FD1S3AX quad_buffer_i7 (.D(quad_count[7]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i7.GSR = "DISABLED";
    FD1S3AX quad_buffer_i6 (.D(quad_count[6]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i6.GSR = "DISABLED";
    FD1S3AX quad_buffer_i5 (.D(quad_count[5]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i5.GSR = "DISABLED";
    FD1S3AX quad_buffer_i4 (.D(quad_count[4]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i4.GSR = "DISABLED";
    FD1S3AX quad_buffer_i3 (.D(quad_count[3]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i3.GSR = "DISABLED";
    FD1S3AX quad_buffer_i2 (.D(quad_count[2]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i2.GSR = "DISABLED";
    FD1S3AX quad_buffer_i1 (.D(quad_count[1]), .CK(\pin_intrpt[8] ), .Q(quad_buffer[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_1553[31] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i31 (.D(\spi_data_out_r_39__N_1553[30] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i30 (.D(\spi_data_out_r_39__N_1553[29] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i29 (.D(\spi_data_out_r_39__N_1553[28] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i28 (.D(\spi_data_out_r_39__N_1553[27] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i27 (.D(\spi_data_out_r_39__N_1553[26] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i26 (.D(\spi_data_out_r_39__N_1553[25] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i25 (.D(\spi_data_out_r_39__N_1553[24] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i24 (.D(\spi_data_out_r_39__N_1553[23] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i23 (.D(\spi_data_out_r_39__N_1553[22] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i22 (.D(\spi_data_out_r_39__N_1553[21] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i21 (.D(\spi_data_out_r_39__N_1553[20] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i20 (.D(\spi_data_out_r_39__N_1553[19] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i19 (.D(\spi_data_out_r_39__N_1553[18] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i18 (.D(\spi_data_out_r_39__N_1553[17] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i17 (.D(\spi_data_out_r_39__N_1553[16] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i16 (.D(\spi_data_out_r_39__N_1553[15] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_1553[14] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_1553[13] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_1553[12] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_1553[11] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_1553[10] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_1553[9] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_1553[8] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_1553[7] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_1553[6] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_1553[5] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_1553[4] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_1553[3] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_1553[2] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_1553[1] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1404[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i2 (.D(quad_b_delayed[1]), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i2.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i1 (.D(quad_b_delayed[0]), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i1.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i31 (.D(n8648), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i31.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i30 (.D(n8650), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i30.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i29 (.D(n8652), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i29.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i28 (.D(n8654), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i28.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i27 (.D(n8656), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i27.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i26 (.D(n8658), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i26.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i25 (.D(n8660), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i25.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i24 (.D(n8662), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i24.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i23 (.D(n8664), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i23.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i22 (.D(n8666), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i22.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i21 (.D(n8668), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i21.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i20 (.D(n8670), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i20.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i19 (.D(n8672), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i19.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i18 (.D(n8674), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i18.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i17 (.D(n8676), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i17.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i16 (.D(n8678), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i16.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i15 (.D(n8680), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i15.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i14 (.D(n8682), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i14.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i13 (.D(n8684), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i13.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i12 (.D(n8686), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i12.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i11 (.D(n8688), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i11.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i10 (.D(n8690), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i10.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i9 (.D(n8692), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i9.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i8 (.D(n8694), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i8.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i7 (.D(n8696), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i7.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i6 (.D(n8698), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i6.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i5 (.D(n8700), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i5.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i4 (.D(n8702), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i4.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i3 (.D(n8704), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i3.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i2 (.D(n8706), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i1 (.D(n8708), .SP(clk_enable_485), .CK(clk), 
            .Q(quad_count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i1.GSR = "DISABLED";
    CCU2D add_1365_7 (.A0(quad_count[4]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[5]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22092), .COUT(n22093), .S0(n4063[4]), .S1(n4063[5]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_7.INIT0 = 16'h5569;
    defparam add_1365_7.INIT1 = 16'h5569;
    defparam add_1365_7.INJECT1_0 = "NO";
    defparam add_1365_7.INJECT1_1 = "NO";
    FD1P3IX quad_homing__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_488), .CD(n30185), 
            .CK(clk), .Q(quad_homing[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(62[8] 69[4])
    defparam quad_homing__i1.GSR = "DISABLED";
    CCU2D add_1365_5 (.A0(quad_count[2]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[3]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22091), .COUT(n22092), .S0(n4063[2]), .S1(n4063[3]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_5.INIT0 = 16'h5569;
    defparam add_1365_5.INIT1 = 16'h5569;
    defparam add_1365_5.INJECT1_0 = "NO";
    defparam add_1365_5.INJECT1_1 = "NO";
    LUT4 i24196_2_lut (.A(resetn_c), .B(quad_homing[1]), .Z(clk_enable_485)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i24196_2_lut.init = 16'h7777;
    LUT4 i3657_4_lut (.A(n4063[0]), .B(quad_set[0]), .C(n5703), .D(n1), 
         .Z(n7981)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i3657_4_lut.init = 16'hc0ca;
    LUT4 i1_4_lut (.A(quad_homing[0]), .B(quad_homing[1]), .C(quad_set_valid), 
         .D(resetn_c), .Z(n5703)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut.init = 16'h1000;
    LUT4 i4324_4_lut (.A(n4063[31]), .B(quad_set[31]), .C(n5703), .D(n1), 
         .Z(n8648)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4324_4_lut.init = 16'hc0ca;
    LUT4 i4326_4_lut (.A(n4063[30]), .B(quad_set[30]), .C(n5703), .D(n1), 
         .Z(n8650)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4326_4_lut.init = 16'hc0ca;
    LUT4 i4328_4_lut (.A(n4063[29]), .B(quad_set[29]), .C(n5703), .D(n1), 
         .Z(n8652)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4328_4_lut.init = 16'hc0ca;
    LUT4 i4330_4_lut (.A(n4063[28]), .B(quad_set[28]), .C(n5703), .D(n1), 
         .Z(n8654)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4330_4_lut.init = 16'hc0ca;
    LUT4 i4332_4_lut (.A(n4063[27]), .B(quad_set[27]), .C(n5703), .D(n1), 
         .Z(n8656)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4332_4_lut.init = 16'hc0ca;
    LUT4 i4334_4_lut (.A(n4063[26]), .B(quad_set[26]), .C(n5703), .D(n1), 
         .Z(n8658)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4334_4_lut.init = 16'hc0ca;
    LUT4 i4336_4_lut (.A(n4063[25]), .B(quad_set[25]), .C(n5703), .D(n1), 
         .Z(n8660)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4336_4_lut.init = 16'hc0ca;
    LUT4 i4338_4_lut (.A(n4063[24]), .B(quad_set[24]), .C(n5703), .D(n1), 
         .Z(n8662)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4338_4_lut.init = 16'hc0ca;
    LUT4 i4340_4_lut (.A(n4063[23]), .B(quad_set[23]), .C(n5703), .D(n1), 
         .Z(n8664)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4340_4_lut.init = 16'hc0ca;
    LUT4 i4342_4_lut (.A(n4063[22]), .B(quad_set[22]), .C(n5703), .D(n1), 
         .Z(n8666)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4342_4_lut.init = 16'hc0ca;
    LUT4 i4344_4_lut (.A(n4063[21]), .B(quad_set[21]), .C(n5703), .D(n1), 
         .Z(n8668)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4344_4_lut.init = 16'hc0ca;
    LUT4 i4346_4_lut (.A(n4063[20]), .B(quad_set[20]), .C(n5703), .D(n1), 
         .Z(n8670)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4346_4_lut.init = 16'hc0ca;
    LUT4 i4348_4_lut (.A(n4063[19]), .B(quad_set[19]), .C(n5703), .D(n1), 
         .Z(n8672)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4348_4_lut.init = 16'hc0ca;
    LUT4 i4350_4_lut (.A(n4063[18]), .B(quad_set[18]), .C(n5703), .D(n1), 
         .Z(n8674)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4350_4_lut.init = 16'hc0ca;
    LUT4 i4352_4_lut (.A(n4063[17]), .B(quad_set[17]), .C(n5703), .D(n1), 
         .Z(n8676)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4352_4_lut.init = 16'hc0ca;
    CCU2D add_1365_3 (.A0(quad_count[0]), .B0(count_dir), .C0(n6), .D0(count_dir), 
          .A1(quad_count[1]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n22090), .COUT(n22091), .S0(n4063[0]), .S1(n4063[1]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_3.INIT0 = 16'h5665;
    defparam add_1365_3.INIT1 = 16'h5569;
    defparam add_1365_3.INJECT1_0 = "NO";
    defparam add_1365_3.INJECT1_1 = "NO";
    LUT4 i4354_4_lut (.A(n4063[16]), .B(quad_set[16]), .C(n5703), .D(n1), 
         .Z(n8678)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4354_4_lut.init = 16'hc0ca;
    LUT4 i4356_4_lut (.A(n4063[15]), .B(quad_set[15]), .C(n5703), .D(n1), 
         .Z(n8680)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4356_4_lut.init = 16'hc0ca;
    LUT4 i4358_4_lut (.A(n4063[14]), .B(quad_set[14]), .C(n5703), .D(n1), 
         .Z(n8682)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4358_4_lut.init = 16'hc0ca;
    LUT4 i4360_4_lut (.A(n4063[13]), .B(quad_set[13]), .C(n5703), .D(n1), 
         .Z(n8684)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4360_4_lut.init = 16'hc0ca;
    LUT4 i4362_4_lut (.A(n4063[12]), .B(quad_set[12]), .C(n5703), .D(n1), 
         .Z(n8686)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4362_4_lut.init = 16'hc0ca;
    CCU2D add_1365_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quad_a_delayed[2]), .B1(quad_b_delayed[1]), .C1(quad_b_delayed[2]), 
          .D1(quad_a_delayed[1]), .COUT(n22090));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1365_1.INIT0 = 16'hF000;
    defparam add_1365_1.INIT1 = 16'h0990;
    defparam add_1365_1.INJECT1_0 = "NO";
    defparam add_1365_1.INJECT1_1 = "NO";
    LUT4 i4364_4_lut (.A(n4063[11]), .B(quad_set[11]), .C(n5703), .D(n1), 
         .Z(n8688)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4364_4_lut.init = 16'hc0ca;
    LUT4 i4366_4_lut (.A(n4063[10]), .B(quad_set[10]), .C(n5703), .D(n1), 
         .Z(n8690)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4366_4_lut.init = 16'hc0ca;
    FD1S3IX quad_a_delayed__i1 (.D(quad_a_delayed[0]), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i1.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i2 (.D(quad_a_delayed[1]), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i2.GSR = "DISABLED";
    LUT4 i4368_4_lut (.A(n4063[9]), .B(quad_set[9]), .C(n5703), .D(n1), 
         .Z(n8692)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4368_4_lut.init = 16'hc0ca;
    LUT4 i4370_4_lut (.A(n4063[8]), .B(quad_set[8]), .C(n5703), .D(n1), 
         .Z(n8694)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4370_4_lut.init = 16'hc0ca;
    LUT4 i4372_4_lut (.A(n4063[7]), .B(quad_set[7]), .C(n5703), .D(n1), 
         .Z(n8696)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4372_4_lut.init = 16'hc0ca;
    LUT4 i4374_4_lut (.A(n4063[6]), .B(quad_set[6]), .C(n5703), .D(n1), 
         .Z(n8698)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4374_4_lut.init = 16'hc0ca;
    LUT4 i4376_4_lut (.A(n4063[5]), .B(quad_set[5]), .C(n5703), .D(n1), 
         .Z(n8700)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4376_4_lut.init = 16'hc0ca;
    LUT4 i4378_4_lut (.A(n4063[4]), .B(quad_set[4]), .C(n5703), .D(n1), 
         .Z(n8702)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4378_4_lut.init = 16'hc0ca;
    LUT4 i4380_4_lut (.A(n4063[3]), .B(quad_set[3]), .C(n5703), .D(n1), 
         .Z(n8704)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4380_4_lut.init = 16'hc0ca;
    LUT4 i4382_4_lut (.A(n4063[2]), .B(quad_set[2]), .C(n5703), .D(n1), 
         .Z(n8706)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4382_4_lut.init = 16'hc0ca;
    LUT4 i4384_4_lut (.A(n4063[1]), .B(quad_set[1]), .C(n5703), .D(n1), 
         .Z(n8708)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4384_4_lut.init = 16'hc0ca;
    LUT4 i2_2_lut (.A(quad_b_delayed[1]), .B(quad_a_delayed[2]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(96[19:96])
    defparam i2_2_lut.init = 16'h6666;
    LUT4 i1_2_lut (.A(quad_a_delayed[1]), .B(quad_b_delayed[2]), .Z(count_dir)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(96[19:96])
    defparam i1_2_lut.init = 16'h6666;
    
endmodule
//
// Verilog Description of module quad_decoder
//

module quad_decoder (quad_count, clk, n30185, \quad_b[0] , \spi_data_out_r_39__N_934[0] , 
            \spi_data_out_r_39__N_1083[0] , quad_buffer, \pin_intrpt[2] , 
            quad_set_valid_N_1158, \quad_a[0] , quad_homing, clk_enable_757, 
            \spi_data_r[0] , clk_enable_807, GND_net, spi_data_out_r_39__N_974, 
            spi_data_out_r_39__N_1163, \spi_cmd_r[2] , \spi_addr_r[7] , 
            n28328, \spi_data_out_r_39__N_934[31] , \spi_data_out_r_39__N_1083[31] , 
            \spi_data_out_r_39__N_934[30] , \spi_data_out_r_39__N_1083[30] , 
            \spi_data_out_r_39__N_934[29] , \spi_data_out_r_39__N_1083[29] , 
            \spi_data_out_r_39__N_934[28] , \spi_data_out_r_39__N_1083[28] , 
            \spi_data_out_r_39__N_934[27] , \spi_data_out_r_39__N_1083[27] , 
            \spi_data_out_r_39__N_934[26] , \spi_data_out_r_39__N_1083[26] , 
            \spi_data_out_r_39__N_934[25] , \spi_data_out_r_39__N_1083[25] , 
            \spi_data_out_r_39__N_934[24] , \spi_data_out_r_39__N_1083[24] , 
            \spi_data_out_r_39__N_934[23] , \spi_data_out_r_39__N_1083[23] , 
            \spi_data_out_r_39__N_934[22] , \spi_data_out_r_39__N_1083[22] , 
            \spi_data_out_r_39__N_934[21] , \spi_data_out_r_39__N_1083[21] , 
            \spi_data_out_r_39__N_934[20] , \spi_data_out_r_39__N_1083[20] , 
            \spi_data_out_r_39__N_934[19] , \spi_data_out_r_39__N_1083[19] , 
            \spi_data_out_r_39__N_934[18] , \spi_data_out_r_39__N_1083[18] , 
            \spi_data_out_r_39__N_934[17] , \spi_data_out_r_39__N_1083[17] , 
            \spi_data_out_r_39__N_934[16] , \spi_data_out_r_39__N_1083[16] , 
            \spi_data_out_r_39__N_934[15] , \spi_data_out_r_39__N_1083[15] , 
            \spi_data_out_r_39__N_934[14] , \spi_data_out_r_39__N_1083[14] , 
            \spi_data_out_r_39__N_934[13] , \spi_data_out_r_39__N_1083[13] , 
            \spi_data_out_r_39__N_934[12] , \spi_data_out_r_39__N_1083[12] , 
            \spi_data_out_r_39__N_934[11] , \spi_data_out_r_39__N_1083[11] , 
            \spi_data_out_r_39__N_934[10] , \spi_data_out_r_39__N_1083[10] , 
            \spi_data_out_r_39__N_934[9] , \spi_data_out_r_39__N_1083[9] , 
            \spi_data_out_r_39__N_934[8] , \spi_data_out_r_39__N_1083[8] , 
            \spi_data_out_r_39__N_934[7] , \spi_data_out_r_39__N_1083[7] , 
            \spi_data_out_r_39__N_934[6] , \spi_data_out_r_39__N_1083[6] , 
            \spi_data_out_r_39__N_934[5] , \spi_data_out_r_39__N_1083[5] , 
            \spi_data_out_r_39__N_934[4] , \spi_data_out_r_39__N_1083[4] , 
            \spi_data_out_r_39__N_934[3] , \spi_data_out_r_39__N_1083[3] , 
            \spi_data_out_r_39__N_934[2] , \spi_data_out_r_39__N_1083[2] , 
            \spi_data_out_r_39__N_934[1] , \spi_data_out_r_39__N_1083[1] , 
            \spi_data_r[1] , \spi_data_r[2] , \spi_data_r[3] , \spi_data_r[4] , 
            \spi_data_r[5] , \spi_data_r[6] , \spi_data_r[7] , \spi_data_r[8] , 
            \spi_data_r[9] , \spi_data_r[10] , \spi_data_r[11] , \spi_data_r[12] , 
            \spi_data_r[13] , \spi_data_r[14] , \spi_data_r[15] , \spi_data_r[16] , 
            \spi_data_r[17] , \spi_data_r[18] , \spi_data_r[19] , \spi_data_r[20] , 
            \spi_data_r[21] , \spi_data_r[22] , \spi_data_r[23] , \spi_data_r[24] , 
            \spi_data_r[25] , \spi_data_r[26] , \spi_data_r[27] , \spi_data_r[28] , 
            \spi_data_r[29] , \spi_data_r[30] , \spi_data_r[31] , n28340, 
            n23916, n26327, quad_set_valid_N_2098, \spi_addr_r[6] , 
            n30209, n28384, \spi_addr_r[2] , n28524, n24169, \spi_addr_r[0] , 
            \spi_addr_r[1] , reset_r_N_4129, n1, resetn_c, n25547) /* synthesis syn_module_defined=1 */ ;
    output [31:0]quad_count;
    input clk;
    input n30185;
    input \quad_b[0] ;
    output \spi_data_out_r_39__N_934[0] ;
    input \spi_data_out_r_39__N_1083[0] ;
    output [31:0]quad_buffer;
    input \pin_intrpt[2] ;
    input quad_set_valid_N_1158;
    input \quad_a[0] ;
    output [1:0]quad_homing;
    input clk_enable_757;
    input \spi_data_r[0] ;
    input clk_enable_807;
    input GND_net;
    output spi_data_out_r_39__N_974;
    input spi_data_out_r_39__N_1163;
    input \spi_cmd_r[2] ;
    input \spi_addr_r[7] ;
    output n28328;
    output \spi_data_out_r_39__N_934[31] ;
    input \spi_data_out_r_39__N_1083[31] ;
    output \spi_data_out_r_39__N_934[30] ;
    input \spi_data_out_r_39__N_1083[30] ;
    output \spi_data_out_r_39__N_934[29] ;
    input \spi_data_out_r_39__N_1083[29] ;
    output \spi_data_out_r_39__N_934[28] ;
    input \spi_data_out_r_39__N_1083[28] ;
    output \spi_data_out_r_39__N_934[27] ;
    input \spi_data_out_r_39__N_1083[27] ;
    output \spi_data_out_r_39__N_934[26] ;
    input \spi_data_out_r_39__N_1083[26] ;
    output \spi_data_out_r_39__N_934[25] ;
    input \spi_data_out_r_39__N_1083[25] ;
    output \spi_data_out_r_39__N_934[24] ;
    input \spi_data_out_r_39__N_1083[24] ;
    output \spi_data_out_r_39__N_934[23] ;
    input \spi_data_out_r_39__N_1083[23] ;
    output \spi_data_out_r_39__N_934[22] ;
    input \spi_data_out_r_39__N_1083[22] ;
    output \spi_data_out_r_39__N_934[21] ;
    input \spi_data_out_r_39__N_1083[21] ;
    output \spi_data_out_r_39__N_934[20] ;
    input \spi_data_out_r_39__N_1083[20] ;
    output \spi_data_out_r_39__N_934[19] ;
    input \spi_data_out_r_39__N_1083[19] ;
    output \spi_data_out_r_39__N_934[18] ;
    input \spi_data_out_r_39__N_1083[18] ;
    output \spi_data_out_r_39__N_934[17] ;
    input \spi_data_out_r_39__N_1083[17] ;
    output \spi_data_out_r_39__N_934[16] ;
    input \spi_data_out_r_39__N_1083[16] ;
    output \spi_data_out_r_39__N_934[15] ;
    input \spi_data_out_r_39__N_1083[15] ;
    output \spi_data_out_r_39__N_934[14] ;
    input \spi_data_out_r_39__N_1083[14] ;
    output \spi_data_out_r_39__N_934[13] ;
    input \spi_data_out_r_39__N_1083[13] ;
    output \spi_data_out_r_39__N_934[12] ;
    input \spi_data_out_r_39__N_1083[12] ;
    output \spi_data_out_r_39__N_934[11] ;
    input \spi_data_out_r_39__N_1083[11] ;
    output \spi_data_out_r_39__N_934[10] ;
    input \spi_data_out_r_39__N_1083[10] ;
    output \spi_data_out_r_39__N_934[9] ;
    input \spi_data_out_r_39__N_1083[9] ;
    output \spi_data_out_r_39__N_934[8] ;
    input \spi_data_out_r_39__N_1083[8] ;
    output \spi_data_out_r_39__N_934[7] ;
    input \spi_data_out_r_39__N_1083[7] ;
    output \spi_data_out_r_39__N_934[6] ;
    input \spi_data_out_r_39__N_1083[6] ;
    output \spi_data_out_r_39__N_934[5] ;
    input \spi_data_out_r_39__N_1083[5] ;
    output \spi_data_out_r_39__N_934[4] ;
    input \spi_data_out_r_39__N_1083[4] ;
    output \spi_data_out_r_39__N_934[3] ;
    input \spi_data_out_r_39__N_1083[3] ;
    output \spi_data_out_r_39__N_934[2] ;
    input \spi_data_out_r_39__N_1083[2] ;
    output \spi_data_out_r_39__N_934[1] ;
    input \spi_data_out_r_39__N_1083[1] ;
    input \spi_data_r[1] ;
    input \spi_data_r[2] ;
    input \spi_data_r[3] ;
    input \spi_data_r[4] ;
    input \spi_data_r[5] ;
    input \spi_data_r[6] ;
    input \spi_data_r[7] ;
    input \spi_data_r[8] ;
    input \spi_data_r[9] ;
    input \spi_data_r[10] ;
    input \spi_data_r[11] ;
    input \spi_data_r[12] ;
    input \spi_data_r[13] ;
    input \spi_data_r[14] ;
    input \spi_data_r[15] ;
    input \spi_data_r[16] ;
    input \spi_data_r[17] ;
    input \spi_data_r[18] ;
    input \spi_data_r[19] ;
    input \spi_data_r[20] ;
    input \spi_data_r[21] ;
    input \spi_data_r[22] ;
    input \spi_data_r[23] ;
    input \spi_data_r[24] ;
    input \spi_data_r[25] ;
    input \spi_data_r[26] ;
    input \spi_data_r[27] ;
    input \spi_data_r[28] ;
    input \spi_data_r[29] ;
    input \spi_data_r[30] ;
    input \spi_data_r[31] ;
    input n28340;
    input n23916;
    input n26327;
    output quad_set_valid_N_2098;
    input \spi_addr_r[6] ;
    input n30209;
    input n28384;
    input \spi_addr_r[2] ;
    input n28524;
    input n24169;
    input \spi_addr_r[0] ;
    input \spi_addr_r[1] ;
    output reset_r_N_4129;
    input n1;
    input resetn_c;
    output n25547;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire \pin_intrpt[2]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[2] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    
    wire n21870, count_dir, n6;
    wire [2:0]quad_b_delayed;   // c:/s_links/sources/quad_decoder.v(35[19:33])
    wire [2:0]quad_a_delayed;   // c:/s_links/sources/quad_decoder.v(34[20:34])
    wire [31:0]n4196;
    
    wire n21871, clk_enable_551, n8552, quad_set_valid;
    wire [31:0]quad_set;   // c:/s_links/sources/quad_decoder.v(39[31:39])
    
    wire n9759, n9757, n9755, n9753, n9751, n9749, n9747, n9745, 
        n9743, n9741, n9739, n9737, n9735, n9733, n9731, n9729, 
        n9727, n9725, n9723, n9721, n9719, n9717, n9715, n9713, 
        n9711, n9709, n9707, n9705, n9703, n9701, n9699, n26325, 
        n5719, n21885, n21884, n21883, n21882, n21881, n21880, 
        n21879, n21878, n21877, n21876, n21875, n21874, n21873, 
        n21872;
    
    CCU2D add_1381_3 (.A0(quad_count[0]), .B0(count_dir), .C0(n6), .D0(count_dir), 
          .A1(quad_count[1]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21870), .COUT(n21871), .S0(n4196[0]), .S1(n4196[1]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_3.INIT0 = 16'h5665;
    defparam add_1381_3.INIT1 = 16'h5569;
    defparam add_1381_3.INJECT1_0 = "NO";
    defparam add_1381_3.INJECT1_1 = "NO";
    FD1P3AX quad_count_i0_i0 (.D(n8552), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i0.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i0 (.D(\quad_b[0] ), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_1083[0] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX quad_buffer_i0 (.D(quad_count[0]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i0.GSR = "DISABLED";
    FD1S3IX quad_set_valid_388 (.D(quad_set_valid_N_1158), .CK(clk), .CD(n30185), 
            .Q(quad_set_valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set_valid_388.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i0 (.D(\quad_a[0] ), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i0.GSR = "DISABLED";
    FD1P3IX quad_homing__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_757), .CD(n30185), 
            .CK(clk), .Q(quad_homing[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(62[8] 69[4])
    defparam quad_homing__i0.GSR = "DISABLED";
    FD1P3IX quad_set__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i0.GSR = "DISABLED";
    CCU2D add_1381_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quad_a_delayed[2]), .B1(quad_b_delayed[1]), .C1(quad_b_delayed[2]), 
          .D1(quad_a_delayed[1]), .COUT(n21870));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_1.INIT0 = 16'hF000;
    defparam add_1381_1.INIT1 = 16'h0990;
    defparam add_1381_1.INJECT1_0 = "NO";
    defparam add_1381_1.INJECT1_1 = "NO";
    FD1S3IX i39_391 (.D(spi_data_out_r_39__N_1163), .CK(clk), .CD(n30185), 
            .Q(spi_data_out_r_39__N_974)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam i39_391.GSR = "DISABLED";
    LUT4 i23626_2_lut (.A(\spi_cmd_r[2] ), .B(\spi_addr_r[7] ), .Z(n28328)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23626_2_lut.init = 16'heeee;
    FD1S3AX quad_buffer_i31 (.D(quad_count[31]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i31.GSR = "DISABLED";
    FD1S3AX quad_buffer_i30 (.D(quad_count[30]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i30.GSR = "DISABLED";
    FD1S3AX quad_buffer_i29 (.D(quad_count[29]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i29.GSR = "DISABLED";
    FD1S3AX quad_buffer_i28 (.D(quad_count[28]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i28.GSR = "DISABLED";
    FD1S3AX quad_buffer_i27 (.D(quad_count[27]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i27.GSR = "DISABLED";
    FD1S3AX quad_buffer_i26 (.D(quad_count[26]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i26.GSR = "DISABLED";
    FD1S3AX quad_buffer_i25 (.D(quad_count[25]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i25.GSR = "DISABLED";
    FD1S3AX quad_buffer_i24 (.D(quad_count[24]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i24.GSR = "DISABLED";
    FD1S3AX quad_buffer_i23 (.D(quad_count[23]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i23.GSR = "DISABLED";
    FD1S3AX quad_buffer_i22 (.D(quad_count[22]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i22.GSR = "DISABLED";
    FD1S3AX quad_buffer_i21 (.D(quad_count[21]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i21.GSR = "DISABLED";
    FD1S3AX quad_buffer_i20 (.D(quad_count[20]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i20.GSR = "DISABLED";
    FD1S3AX quad_buffer_i19 (.D(quad_count[19]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i19.GSR = "DISABLED";
    FD1S3AX quad_buffer_i18 (.D(quad_count[18]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i18.GSR = "DISABLED";
    FD1S3AX quad_buffer_i17 (.D(quad_count[17]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i17.GSR = "DISABLED";
    FD1S3AX quad_buffer_i16 (.D(quad_count[16]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i16.GSR = "DISABLED";
    FD1S3AX quad_buffer_i15 (.D(quad_count[15]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i15.GSR = "DISABLED";
    FD1S3AX quad_buffer_i14 (.D(quad_count[14]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i14.GSR = "DISABLED";
    FD1S3AX quad_buffer_i13 (.D(quad_count[13]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i13.GSR = "DISABLED";
    FD1S3AX quad_buffer_i12 (.D(quad_count[12]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i12.GSR = "DISABLED";
    FD1S3AX quad_buffer_i11 (.D(quad_count[11]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i11.GSR = "DISABLED";
    FD1S3AX quad_buffer_i10 (.D(quad_count[10]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i10.GSR = "DISABLED";
    FD1S3AX quad_buffer_i9 (.D(quad_count[9]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i9.GSR = "DISABLED";
    FD1S3AX quad_buffer_i8 (.D(quad_count[8]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i8.GSR = "DISABLED";
    FD1S3AX quad_buffer_i7 (.D(quad_count[7]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i7.GSR = "DISABLED";
    FD1S3AX quad_buffer_i6 (.D(quad_count[6]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i6.GSR = "DISABLED";
    FD1S3AX quad_buffer_i5 (.D(quad_count[5]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i5.GSR = "DISABLED";
    FD1S3AX quad_buffer_i4 (.D(quad_count[4]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i4.GSR = "DISABLED";
    FD1S3AX quad_buffer_i3 (.D(quad_count[3]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i3.GSR = "DISABLED";
    FD1S3AX quad_buffer_i2 (.D(quad_count[2]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i2.GSR = "DISABLED";
    FD1S3AX quad_buffer_i1 (.D(quad_count[1]), .CK(\pin_intrpt[2] ), .Q(quad_buffer[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(139[8] 141[4])
    defparam quad_buffer_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_1083[31] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i31 (.D(\spi_data_out_r_39__N_1083[30] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i30 (.D(\spi_data_out_r_39__N_1083[29] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i29 (.D(\spi_data_out_r_39__N_1083[28] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i28 (.D(\spi_data_out_r_39__N_1083[27] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i27 (.D(\spi_data_out_r_39__N_1083[26] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i26 (.D(\spi_data_out_r_39__N_1083[25] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i25 (.D(\spi_data_out_r_39__N_1083[24] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i24 (.D(\spi_data_out_r_39__N_1083[23] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i23 (.D(\spi_data_out_r_39__N_1083[22] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i22 (.D(\spi_data_out_r_39__N_1083[21] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i21 (.D(\spi_data_out_r_39__N_1083[20] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i20 (.D(\spi_data_out_r_39__N_1083[19] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i19 (.D(\spi_data_out_r_39__N_1083[18] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i18 (.D(\spi_data_out_r_39__N_1083[17] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i17 (.D(\spi_data_out_r_39__N_1083[16] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i16 (.D(\spi_data_out_r_39__N_1083[15] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_1083[14] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_1083[13] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_1083[12] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_1083[11] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_1083[10] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_1083[9] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_1083[8] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_1083[7] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_1083[6] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_1083[5] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_1083[4] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_1083[3] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_1083[2] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_1083[1] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(72[8] 81[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i2 (.D(quad_b_delayed[1]), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i2.GSR = "DISABLED";
    FD1S3IX quad_b_delayed__i1 (.D(quad_b_delayed[0]), .CK(clk), .CD(n30185), 
            .Q(quad_b_delayed[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_b_delayed__i1.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i31 (.D(n9759), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i31.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i30 (.D(n9757), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i30.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i29 (.D(n9755), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i29.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i28 (.D(n9753), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i28.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i27 (.D(n9751), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i27.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i26 (.D(n9749), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i26.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i25 (.D(n9747), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i25.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i24 (.D(n9745), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i24.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i23 (.D(n9743), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i23.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i22 (.D(n9741), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i22.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i21 (.D(n9739), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i21.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i20 (.D(n9737), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i20.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i19 (.D(n9735), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i19.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i18 (.D(n9733), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i18.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i17 (.D(n9731), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i17.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i16 (.D(n9729), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i16.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i15 (.D(n9727), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i15.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i14 (.D(n9725), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i14.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i13 (.D(n9723), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i13.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i12 (.D(n9721), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i12.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i11 (.D(n9719), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i11.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i10 (.D(n9717), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i10.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i9 (.D(n9715), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i9.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i8 (.D(n9713), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i8.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i7 (.D(n9711), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i7.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i6 (.D(n9709), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i6.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i5 (.D(n9707), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i5.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i4 (.D(n9705), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i4.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i3 (.D(n9703), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i3.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i2 (.D(n9701), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i1 (.D(n9699), .SP(clk_enable_551), .CK(clk), 
            .Q(quad_count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(100[8] 137[4])
    defparam quad_count_i0_i1.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i1 (.D(quad_a_delayed[0]), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i1.GSR = "DISABLED";
    FD1S3IX quad_a_delayed__i2 (.D(quad_a_delayed[1]), .CK(clk), .CD(n30185), 
            .Q(quad_a_delayed[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(85[8] 94[4])
    defparam quad_a_delayed__i2.GSR = "DISABLED";
    FD1P3IX quad_homing__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_757), .CD(n30185), 
            .CK(clk), .Q(quad_homing[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(62[8] 69[4])
    defparam quad_homing__i1.GSR = "DISABLED";
    FD1P3IX quad_set__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i1.GSR = "DISABLED";
    FD1P3IX quad_set__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i2.GSR = "DISABLED";
    FD1P3IX quad_set__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i3.GSR = "DISABLED";
    FD1P3IX quad_set__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i4.GSR = "DISABLED";
    FD1P3IX quad_set__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i5.GSR = "DISABLED";
    FD1P3IX quad_set__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i6.GSR = "DISABLED";
    FD1P3IX quad_set__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i7.GSR = "DISABLED";
    FD1P3IX quad_set__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i8.GSR = "DISABLED";
    FD1P3IX quad_set__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i9.GSR = "DISABLED";
    FD1P3IX quad_set__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i10.GSR = "DISABLED";
    FD1P3IX quad_set__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i11.GSR = "DISABLED";
    FD1P3IX quad_set__i12 (.D(\spi_data_r[12] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i12.GSR = "DISABLED";
    FD1P3IX quad_set__i13 (.D(\spi_data_r[13] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i13.GSR = "DISABLED";
    FD1P3IX quad_set__i14 (.D(\spi_data_r[14] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i14.GSR = "DISABLED";
    FD1P3IX quad_set__i15 (.D(\spi_data_r[15] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i15.GSR = "DISABLED";
    FD1P3IX quad_set__i16 (.D(\spi_data_r[16] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i16.GSR = "DISABLED";
    FD1P3IX quad_set__i17 (.D(\spi_data_r[17] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i17.GSR = "DISABLED";
    FD1P3IX quad_set__i18 (.D(\spi_data_r[18] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i18.GSR = "DISABLED";
    FD1P3IX quad_set__i19 (.D(\spi_data_r[19] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i19.GSR = "DISABLED";
    FD1P3IX quad_set__i20 (.D(\spi_data_r[20] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i20.GSR = "DISABLED";
    FD1P3IX quad_set__i21 (.D(\spi_data_r[21] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i21.GSR = "DISABLED";
    FD1P3IX quad_set__i22 (.D(\spi_data_r[22] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i22.GSR = "DISABLED";
    FD1P3IX quad_set__i23 (.D(\spi_data_r[23] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i23.GSR = "DISABLED";
    FD1P3IX quad_set__i24 (.D(\spi_data_r[24] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i24.GSR = "DISABLED";
    FD1P3IX quad_set__i25 (.D(\spi_data_r[25] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i25.GSR = "DISABLED";
    FD1P3IX quad_set__i26 (.D(\spi_data_r[26] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i26.GSR = "DISABLED";
    FD1P3IX quad_set__i27 (.D(\spi_data_r[27] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i27.GSR = "DISABLED";
    FD1P3IX quad_set__i28 (.D(\spi_data_r[28] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i28.GSR = "DISABLED";
    FD1P3IX quad_set__i29 (.D(\spi_data_r[29] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i29.GSR = "DISABLED";
    FD1P3IX quad_set__i30 (.D(\spi_data_r[30] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i30.GSR = "DISABLED";
    FD1P3IX quad_set__i31 (.D(\spi_data_r[31] ), .SP(clk_enable_807), .CD(n30185), 
            .CK(clk), .Q(quad_set[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=263, LSE_RLINE=283 */ ;   // c:/s_links/sources/quad_decoder.v(47[8] 60[4])
    defparam quad_set__i31.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(n28340), .B(n23916), .C(n26327), .D(n26325), .Z(quad_set_valid_N_2098)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_4_lut.init = 16'h4000;
    LUT4 i1_4_lut_adj_586 (.A(\spi_addr_r[6] ), .B(n30209), .C(n28384), 
         .D(\spi_addr_r[2] ), .Z(n26325)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_586.init = 16'h0100;
    LUT4 i1_4_lut_adj_587 (.A(n28524), .B(n24169), .C(\spi_addr_r[0] ), 
         .D(\spi_addr_r[1] ), .Z(reset_r_N_4129)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_587.init = 16'h0004;
    LUT4 i5435_4_lut (.A(n4196[31]), .B(quad_set[31]), .C(n5719), .D(n1), 
         .Z(n9759)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5435_4_lut.init = 16'hc0ca;
    LUT4 i5433_4_lut (.A(n4196[30]), .B(quad_set[30]), .C(n5719), .D(n1), 
         .Z(n9757)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5433_4_lut.init = 16'hc0ca;
    LUT4 i5431_4_lut (.A(n4196[29]), .B(quad_set[29]), .C(n5719), .D(n1), 
         .Z(n9755)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5431_4_lut.init = 16'hc0ca;
    LUT4 i5429_4_lut (.A(n4196[28]), .B(quad_set[28]), .C(n5719), .D(n1), 
         .Z(n9753)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5429_4_lut.init = 16'hc0ca;
    LUT4 i5427_4_lut (.A(n4196[27]), .B(quad_set[27]), .C(n5719), .D(n1), 
         .Z(n9751)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5427_4_lut.init = 16'hc0ca;
    LUT4 i5425_4_lut (.A(n4196[26]), .B(quad_set[26]), .C(n5719), .D(n1), 
         .Z(n9749)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5425_4_lut.init = 16'hc0ca;
    LUT4 i5423_4_lut (.A(n4196[25]), .B(quad_set[25]), .C(n5719), .D(n1), 
         .Z(n9747)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5423_4_lut.init = 16'hc0ca;
    LUT4 i1_4_lut_adj_588 (.A(\spi_addr_r[7] ), .B(\spi_addr_r[0] ), .C(\spi_addr_r[2] ), 
         .D(resetn_c), .Z(n25547)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_588.init = 16'h0100;
    LUT4 i5421_4_lut (.A(n4196[24]), .B(quad_set[24]), .C(n5719), .D(n1), 
         .Z(n9745)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5421_4_lut.init = 16'hc0ca;
    LUT4 i5419_4_lut (.A(n4196[23]), .B(quad_set[23]), .C(n5719), .D(n1), 
         .Z(n9743)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5419_4_lut.init = 16'hc0ca;
    LUT4 i5417_4_lut (.A(n4196[22]), .B(quad_set[22]), .C(n5719), .D(n1), 
         .Z(n9741)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5417_4_lut.init = 16'hc0ca;
    LUT4 i5415_4_lut (.A(n4196[21]), .B(quad_set[21]), .C(n5719), .D(n1), 
         .Z(n9739)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5415_4_lut.init = 16'hc0ca;
    LUT4 i5413_4_lut (.A(n4196[20]), .B(quad_set[20]), .C(n5719), .D(n1), 
         .Z(n9737)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5413_4_lut.init = 16'hc0ca;
    LUT4 i5411_4_lut (.A(n4196[19]), .B(quad_set[19]), .C(n5719), .D(n1), 
         .Z(n9735)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5411_4_lut.init = 16'hc0ca;
    LUT4 i5409_4_lut (.A(n4196[18]), .B(quad_set[18]), .C(n5719), .D(n1), 
         .Z(n9733)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5409_4_lut.init = 16'hc0ca;
    LUT4 i5407_4_lut (.A(n4196[17]), .B(quad_set[17]), .C(n5719), .D(n1), 
         .Z(n9731)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5407_4_lut.init = 16'hc0ca;
    LUT4 i5405_4_lut (.A(n4196[16]), .B(quad_set[16]), .C(n5719), .D(n1), 
         .Z(n9729)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5405_4_lut.init = 16'hc0ca;
    LUT4 i5403_4_lut (.A(n4196[15]), .B(quad_set[15]), .C(n5719), .D(n1), 
         .Z(n9727)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5403_4_lut.init = 16'hc0ca;
    LUT4 i5401_4_lut (.A(n4196[14]), .B(quad_set[14]), .C(n5719), .D(n1), 
         .Z(n9725)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5401_4_lut.init = 16'hc0ca;
    LUT4 i5399_4_lut (.A(n4196[13]), .B(quad_set[13]), .C(n5719), .D(n1), 
         .Z(n9723)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5399_4_lut.init = 16'hc0ca;
    LUT4 i5397_4_lut (.A(n4196[12]), .B(quad_set[12]), .C(n5719), .D(n1), 
         .Z(n9721)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5397_4_lut.init = 16'hc0ca;
    LUT4 i5395_4_lut (.A(n4196[11]), .B(quad_set[11]), .C(n5719), .D(n1), 
         .Z(n9719)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5395_4_lut.init = 16'hc0ca;
    LUT4 i5393_4_lut (.A(n4196[10]), .B(quad_set[10]), .C(n5719), .D(n1), 
         .Z(n9717)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5393_4_lut.init = 16'hc0ca;
    LUT4 i5391_4_lut (.A(n4196[9]), .B(quad_set[9]), .C(n5719), .D(n1), 
         .Z(n9715)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5391_4_lut.init = 16'hc0ca;
    LUT4 i5389_4_lut (.A(n4196[8]), .B(quad_set[8]), .C(n5719), .D(n1), 
         .Z(n9713)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5389_4_lut.init = 16'hc0ca;
    LUT4 i5387_4_lut (.A(n4196[7]), .B(quad_set[7]), .C(n5719), .D(n1), 
         .Z(n9711)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5387_4_lut.init = 16'hc0ca;
    LUT4 i5385_4_lut (.A(n4196[6]), .B(quad_set[6]), .C(n5719), .D(n1), 
         .Z(n9709)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5385_4_lut.init = 16'hc0ca;
    LUT4 i5383_4_lut (.A(n4196[5]), .B(quad_set[5]), .C(n5719), .D(n1), 
         .Z(n9707)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5383_4_lut.init = 16'hc0ca;
    LUT4 i5381_4_lut (.A(n4196[4]), .B(quad_set[4]), .C(n5719), .D(n1), 
         .Z(n9705)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5381_4_lut.init = 16'hc0ca;
    LUT4 i2_2_lut (.A(quad_b_delayed[1]), .B(quad_a_delayed[2]), .Z(n6)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(96[19:96])
    defparam i2_2_lut.init = 16'h6666;
    LUT4 i5379_4_lut (.A(n4196[3]), .B(quad_set[3]), .C(n5719), .D(n1), 
         .Z(n9703)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5379_4_lut.init = 16'hc0ca;
    LUT4 i5377_4_lut (.A(n4196[2]), .B(quad_set[2]), .C(n5719), .D(n1), 
         .Z(n9701)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5377_4_lut.init = 16'hc0ca;
    LUT4 i5375_4_lut (.A(n4196[1]), .B(quad_set[1]), .C(n5719), .D(n1), 
         .Z(n9699)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i5375_4_lut.init = 16'hc0ca;
    CCU2D add_1381_33 (.A0(quad_count[30]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[31]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21885), .S0(n4196[30]), .S1(n4196[31]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_33.INIT0 = 16'h5569;
    defparam add_1381_33.INIT1 = 16'h5569;
    defparam add_1381_33.INJECT1_0 = "NO";
    defparam add_1381_33.INJECT1_1 = "NO";
    CCU2D add_1381_31 (.A0(quad_count[28]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[29]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21884), .COUT(n21885), .S0(n4196[28]), .S1(n4196[29]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_31.INIT0 = 16'h5569;
    defparam add_1381_31.INIT1 = 16'h5569;
    defparam add_1381_31.INJECT1_0 = "NO";
    defparam add_1381_31.INJECT1_1 = "NO";
    CCU2D add_1381_29 (.A0(quad_count[26]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[27]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21883), .COUT(n21884), .S0(n4196[26]), .S1(n4196[27]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_29.INIT0 = 16'h5569;
    defparam add_1381_29.INIT1 = 16'h5569;
    defparam add_1381_29.INJECT1_0 = "NO";
    defparam add_1381_29.INJECT1_1 = "NO";
    CCU2D add_1381_27 (.A0(quad_count[24]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[25]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21882), .COUT(n21883), .S0(n4196[24]), .S1(n4196[25]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_27.INIT0 = 16'h5569;
    defparam add_1381_27.INIT1 = 16'h5569;
    defparam add_1381_27.INJECT1_0 = "NO";
    defparam add_1381_27.INJECT1_1 = "NO";
    CCU2D add_1381_25 (.A0(quad_count[22]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[23]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21881), .COUT(n21882), .S0(n4196[22]), .S1(n4196[23]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_25.INIT0 = 16'h5569;
    defparam add_1381_25.INIT1 = 16'h5569;
    defparam add_1381_25.INJECT1_0 = "NO";
    defparam add_1381_25.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(quad_a_delayed[1]), .B(quad_b_delayed[2]), .Z(count_dir)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(96[19:96])
    defparam i1_2_lut.init = 16'h6666;
    CCU2D add_1381_23 (.A0(quad_count[20]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[21]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21880), .COUT(n21881), .S0(n4196[20]), .S1(n4196[21]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_23.INIT0 = 16'h5569;
    defparam add_1381_23.INIT1 = 16'h5569;
    defparam add_1381_23.INJECT1_0 = "NO";
    defparam add_1381_23.INJECT1_1 = "NO";
    CCU2D add_1381_21 (.A0(quad_count[18]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[19]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21879), .COUT(n21880), .S0(n4196[18]), .S1(n4196[19]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_21.INIT0 = 16'h5569;
    defparam add_1381_21.INIT1 = 16'h5569;
    defparam add_1381_21.INJECT1_0 = "NO";
    defparam add_1381_21.INJECT1_1 = "NO";
    CCU2D add_1381_19 (.A0(quad_count[16]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[17]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21878), .COUT(n21879), .S0(n4196[16]), .S1(n4196[17]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_19.INIT0 = 16'h5569;
    defparam add_1381_19.INIT1 = 16'h5569;
    defparam add_1381_19.INJECT1_0 = "NO";
    defparam add_1381_19.INJECT1_1 = "NO";
    CCU2D add_1381_17 (.A0(quad_count[14]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[15]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21877), .COUT(n21878), .S0(n4196[14]), .S1(n4196[15]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_17.INIT0 = 16'h5569;
    defparam add_1381_17.INIT1 = 16'h5569;
    defparam add_1381_17.INJECT1_0 = "NO";
    defparam add_1381_17.INJECT1_1 = "NO";
    CCU2D add_1381_15 (.A0(quad_count[12]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[13]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21876), .COUT(n21877), .S0(n4196[12]), .S1(n4196[13]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_15.INIT0 = 16'h5569;
    defparam add_1381_15.INIT1 = 16'h5569;
    defparam add_1381_15.INJECT1_0 = "NO";
    defparam add_1381_15.INJECT1_1 = "NO";
    CCU2D add_1381_13 (.A0(quad_count[10]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[11]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21875), .COUT(n21876), .S0(n4196[10]), .S1(n4196[11]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_13.INIT0 = 16'h5569;
    defparam add_1381_13.INIT1 = 16'h5569;
    defparam add_1381_13.INJECT1_0 = "NO";
    defparam add_1381_13.INJECT1_1 = "NO";
    CCU2D add_1381_11 (.A0(quad_count[8]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[9]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21874), .COUT(n21875), .S0(n4196[8]), .S1(n4196[9]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_11.INIT0 = 16'h5569;
    defparam add_1381_11.INIT1 = 16'h5569;
    defparam add_1381_11.INJECT1_0 = "NO";
    defparam add_1381_11.INJECT1_1 = "NO";
    CCU2D add_1381_9 (.A0(quad_count[6]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[7]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21873), .COUT(n21874), .S0(n4196[6]), .S1(n4196[7]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_9.INIT0 = 16'h5569;
    defparam add_1381_9.INIT1 = 16'h5569;
    defparam add_1381_9.INJECT1_0 = "NO";
    defparam add_1381_9.INJECT1_1 = "NO";
    CCU2D add_1381_7 (.A0(quad_count[4]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[5]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21872), .COUT(n21873), .S0(n4196[4]), .S1(n4196[5]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_7.INIT0 = 16'h5569;
    defparam add_1381_7.INIT1 = 16'h5569;
    defparam add_1381_7.INJECT1_0 = "NO";
    defparam add_1381_7.INJECT1_1 = "NO";
    CCU2D add_1381_5 (.A0(quad_count[2]), .B0(quad_b_delayed[2]), .C0(quad_a_delayed[1]), 
          .D0(n6), .A1(quad_count[3]), .B1(quad_b_delayed[2]), .C1(quad_a_delayed[1]), 
          .D1(n6), .CIN(n21871), .COUT(n21872), .S0(n4196[2]), .S1(n4196[3]));   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam add_1381_5.INIT0 = 16'h5569;
    defparam add_1381_5.INIT1 = 16'h5569;
    defparam add_1381_5.INJECT1_0 = "NO";
    defparam add_1381_5.INJECT1_1 = "NO";
    LUT4 i24205_2_lut (.A(resetn_c), .B(quad_homing[1]), .Z(clk_enable_551)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i24205_2_lut.init = 16'h7777;
    LUT4 i4228_4_lut (.A(n4196[0]), .B(quad_set[0]), .C(n5719), .D(n1), 
         .Z(n8552)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(105[7] 136[5])
    defparam i4228_4_lut.init = 16'hc0ca;
    LUT4 i1_4_lut_adj_589 (.A(quad_homing[0]), .B(quad_homing[1]), .C(quad_set_valid), 
         .D(resetn_c), .Z(n5719)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_589.init = 16'h1000;
    
endmodule
//
// Verilog Description of module \stepper(DEV_ID=6,UART_ADDRESS_WIDTH=4) 
//

module \stepper(DEV_ID=6,UART_ADDRESS_WIDTH=4)  (\spi_data_out_r_39__N_5540[4] , 
            spi_data_out_r_39__N_5580, \spi_data_out_r_39__N_4511[4] , spi_data_out_r_39__N_4551, 
            clk, \spi_data_out_r_39__N_1404[4] , \spi_data_out_r_39__N_1639[4] , 
            spi_data_out_r_39__N_1444, spi_data_out_r_39__N_1679, \spi_data_out_r_39__N_1874[4] , 
            spi_data_out_r_39__N_1914, \spi_data_out_r_39__N_1169[4] , spi_data_out_r_39__N_1209, 
            \spi_data_out_r_39__N_2109[4] , \spi_data_out_r_39__N_934[4] , 
            spi_data_out_r_39__N_2149, spi_data_out_r_39__N_974, \spi_data_out_r_39__N_2344[4] , 
            spi_data_out_r_39__N_2384, \spi_data_out_r_39__N_5197[4] , \spi_data_out_r_39__N_4854[4] , 
            spi_data_out_r_39__N_5237, spi_data_out_r_39__N_4894, spi_data_out_r_39__N_5923, 
            \spi_data_out_r[5] , \spi_data_out_r_39__N_3825[5] , \spi_data_out_r_39__N_4168[5] , 
            spi_data_out_r_39__N_3865, spi_data_out_r_39__N_4208, \spi_data_out_r_39__N_5540[5] , 
            reset_r, n30185, n30028, NSL, clk_1MHz, \spi_data_out_r_39__N_4511[5] , 
            \spi_data_out_r_39__N_1404[5] , \spi_data_out_r_39__N_1639[5] , 
            \spi_data_out_r_39__N_1874[5] , \spi_data_out_r_39__N_1169[5] , 
            \spi_data_out_r_39__N_2109[5] , \spi_data_out_r_39__N_934[5] , 
            \spi_data_out_r_39__N_2344[5] , \spi_data_out_r_39__N_5197[5] , 
            \spi_data_out_r_39__N_4854[5] , clk_enable_180, \spi_data_r[0] , 
            \spi_data_out_r[6] , \spi_data_out_r_39__N_3825[6] , \spi_data_out_r_39__N_4168[6] , 
            \spi_data_out_r_39__N_5540[6] , \spi_data_out_r_39__N_4511[6] , 
            \spi_data_out_r_39__N_1404[6] , \spi_data_out_r_39__N_1639[6] , 
            \spi_data_out_r_39__N_1874[6] , \spi_data_out_r_39__N_1169[6] , 
            \spi_data_out_r_39__N_2109[6] , \spi_data_out_r_39__N_934[6] , 
            \spi_data_out_r_39__N_2344[6] , \spi_data_out_r_39__N_5197[6] , 
            \spi_data_out_r_39__N_4854[6] , \spi_data_out_r[7] , \spi_data_out_r_39__N_3825[7] , 
            \spi_data_out_r_39__N_4168[7] , \spi_data_out_r_39__N_5540[7] , 
            \spi_data_out_r_39__N_4511[7] , \spi_data_out_r_39__N_1404[7] , 
            \spi_data_out_r_39__N_1639[7] , n30143, \spi_data_out_r_39__N_1874[7] , 
            \spi_data_out_r_39__N_1169[7] , \spi_data_out_r_39__N_2109[7] , 
            \spi_data_out_r_39__N_934[7] , \spi_data_out_r_39__N_2344[7] , 
            \spi_data_out_r_39__N_5197[7] , \spi_data_out_r_39__N_4854[7] , 
            resetn_c, \spi_data_out_r[10] , \spi_data_out_r_39__N_3825[10] , 
            \spi_data_out_r_39__N_4168[10] , \spi_data_r[2] , \spi_data_r[1] , 
            \spi_data_out_r_39__N_5540[10] , \spi_data_out_r_39__N_4511[10] , 
            \spi_data_out_r_39__N_1404[10] , \spi_data_out_r_39__N_1639[10] , 
            \spi_data_out_r_39__N_1874[10] , \spi_data_out_r_39__N_1169[10] , 
            \spi_data_out_r_39__N_2109[10] , \spi_data_out_r_39__N_934[10] , 
            \spi_data_out_r_39__N_2344[10] , \spi_data_out_r_39__N_5197[10] , 
            \spi_data_out_r_39__N_4854[10] , \spi_data_out_r[11] , \spi_data_out_r_39__N_3825[11] , 
            \spi_data_out_r_39__N_4168[11] , \spi_data_out_r_39__N_5540[11] , 
            \spi_data_out_r_39__N_4511[11] , \spi_data_out_r_39__N_1404[11] , 
            \spi_data_out_r_39__N_1639[11] , \spi_data_out_r_39__N_1874[11] , 
            \spi_data_out_r_39__N_1169[11] , \spi_data_out_r_39__N_2109[11] , 
            \spi_data_out_r_39__N_934[11] , \spi_data_out_r_39__N_2344[11] , 
            \spi_data_out_r_39__N_5197[11] , \spi_data_out_r_39__N_4854[11] , 
            \spi_data_out_r[12] , \spi_data_out_r_39__N_3825[12] , \spi_data_out_r_39__N_4168[12] , 
            \spi_data_out_r_39__N_5540[12] , \spi_data_out_r_39__N_4511[12] , 
            \spi_data_out_r_39__N_1404[12] , \spi_data_out_r_39__N_1639[12] , 
            \spi_data_out_r_39__N_1874[12] , \spi_data_out_r_39__N_1169[12] , 
            \spi_data_out_r_39__N_2109[12] , \spi_data_out_r_39__N_934[12] , 
            \spi_data_out_r_39__N_2344[12] , \spi_data_out_r_39__N_5197[12] , 
            \spi_data_out_r_39__N_4854[12] , \spi_data_out_r[13] , \spi_data_out_r_39__N_3825[13] , 
            \spi_data_out_r_39__N_4168[13] , digital_output_r, clk_enable_222, 
            n28550, \spi_data_out_r_39__N_5540[13] , EM_STOP, n25741, 
            n23916, \spi_data_out_r_39__N_4511[13] , \spi_data_out_r_39__N_1404[13] , 
            \spi_data_out_r_39__N_1639[13] , \spi_data_out_r_39__N_1874[13] , 
            \spi_data_out_r_39__N_1169[13] , \spi_data_out_r_39__N_2109[13] , 
            \spi_data_out_r_39__N_934[13] , \spi_data_out_r_39__N_2344[13] , 
            \spi_data_out_r_39__N_5197[13] , \spi_data_out_r_39__N_4854[13] , 
            \spi_data_out_r[14] , \spi_data_out_r_39__N_3825[14] , \spi_data_out_r_39__N_4168[14] , 
            \spi_data_out_r_39__N_5540[14] , \spi_data_out_r_39__N_4511[14] , 
            \spi_data_out_r_39__N_1404[14] , \spi_data_out_r_39__N_1639[14] , 
            \spi_data_out_r_39__N_1874[14] , \spi_data_out_r_39__N_1169[14] , 
            \spi_data_out_r_39__N_2109[14] , \spi_data_out_r_39__N_934[14] , 
            \spi_data_out_r_39__N_2344[14] , \spi_data_out_r_39__N_5197[14] , 
            \spi_data_out_r_39__N_4854[14] , \spi_data_out_r[15] , \spi_data_out_r_39__N_3825[15] , 
            \spi_data_out_r_39__N_4168[15] , \spi_data_out_r_39__N_5540[15] , 
            \spi_data_out_r_39__N_4511[15] , \spi_data_out_r_39__N_1404[15] , 
            \spi_data_out_r_39__N_1639[15] , \spi_data_out_r_39__N_1874[15] , 
            \spi_data_out_r_39__N_1169[15] , \spi_data_out_r_39__N_2109[15] , 
            \spi_data_out_r_39__N_934[15] , \spi_data_out_r_39__N_2344[15] , 
            \spi_data_out_r_39__N_5197[15] , \spi_data_out_r_39__N_4854[15] , 
            \spi_data_out_r[16] , \spi_data_out_r_39__N_3825[16] , \spi_data_out_r_39__N_4168[16] , 
            \spi_data_out_r_39__N_5540[16] , \spi_data_out_r_39__N_4511[16] , 
            \spi_data_out_r_39__N_1404[16] , \spi_data_out_r_39__N_1639[16] , 
            \spi_data_out_r_39__N_1874[16] , \spi_data_out_r_39__N_1169[16] , 
            \spi_data_out_r_39__N_2109[16] , \spi_data_out_r_39__N_934[16] , 
            \spi_data_out_r_39__N_2344[16] , \spi_data_out_r_39__N_5197[16] , 
            \spi_data_out_r_39__N_4854[16] , \spi_data_out_r[17] , \spi_data_out_r_39__N_3825[17] , 
            \spi_data_out_r_39__N_4168[17] , \spi_data_out_r_39__N_5540[17] , 
            \spi_data_out_r_39__N_4511[17] , \spi_data_out_r_39__N_1404[17] , 
            \spi_data_out_r_39__N_1639[17] , spi_data_out_r_39__N_6220, 
            \spi_data_out_r_39__N_1874[17] , \spi_data_out_r_39__N_1169[17] , 
            \spi_data_out_r_39__N_2109[17] , \spi_data_out_r_39__N_934[17] , 
            \spi_data_out_r_39__N_2344[17] , \spi_data_out_r_39__N_5197[17] , 
            \spi_data_out_r_39__N_4854[17] , \spi_data_out_r[18] , \spi_data_out_r_39__N_3825[18] , 
            \spi_data_out_r_39__N_4168[18] , \spi_data_out_r_39__N_5540[18] , 
            \spi_data_out_r_39__N_4511[18] , \spi_data_out_r_39__N_1404[18] , 
            \spi_data_out_r_39__N_1639[18] , \spi_data_out_r_39__N_1874[18] , 
            \spi_data_out_r_39__N_1169[18] , \spi_data_out_r_39__N_2109[18] , 
            \spi_data_out_r_39__N_934[18] , \spi_data_out_r_39__N_2344[18] , 
            \spi_data_out_r_39__N_5197[18] , \spi_data_out_r_39__N_4854[18] , 
            \spi_data_out_r[19] , \spi_data_out_r_39__N_3825[19] , \spi_data_out_r_39__N_4168[19] , 
            \spi_data_out_r_39__N_5540[19] , \spi_data_out_r_39__N_4511[19] , 
            \spi_data_out_r_39__N_1404[19] , \spi_data_out_r_39__N_1639[19] , 
            \spi_data_out_r_39__N_1874[19] , \spi_data_out_r_39__N_1169[19] , 
            \spi_data_out_r_39__N_2109[19] , \spi_data_out_r_39__N_934[19] , 
            \spi_data_out_r_39__N_2344[19] , \spi_data_out_r_39__N_5197[19] , 
            \spi_data_out_r_39__N_4854[19] , \spi_data_out_r[20] , \spi_data_out_r_39__N_3825[20] , 
            \spi_data_out_r_39__N_4168[20] , \spi_data_out_r_39__N_5540[20] , 
            \spi_data_out_r_39__N_4511[20] , \spi_data_out_r_39__N_1404[20] , 
            \spi_data_out_r_39__N_1639[20] , \spi_data_out_r_39__N_1874[20] , 
            \spi_data_out_r_39__N_1169[20] , \spi_data_out_r_39__N_2109[20] , 
            \spi_data_out_r_39__N_934[20] , \spi_data_out_r_39__N_2344[20] , 
            \spi_data_out_r_39__N_5197[20] , \spi_data_out_r_39__N_4854[20] , 
            \spi_data_out_r[21] , \spi_data_out_r_39__N_3825[21] , \spi_data_out_r_39__N_4168[21] , 
            \spi_data_out_r_39__N_5540[21] , \spi_data_out_r_39__N_4511[21] , 
            \spi_data_out_r_39__N_1404[21] , \spi_data_out_r_39__N_1639[21] , 
            \spi_data_out_r_39__N_1874[21] , \spi_data_out_r_39__N_1169[21] , 
            \spi_data_out_r_39__N_2109[21] , \spi_data_out_r_39__N_934[21] , 
            \spi_data_out_r_39__N_2344[21] , \spi_data_out_r_39__N_5197[21] , 
            \spi_data_out_r_39__N_4854[21] , \spi_data_out_r[22] , \spi_data_out_r_39__N_3825[22] , 
            \spi_data_out_r_39__N_4168[22] , \spi_data_out_r_39__N_5540[22] , 
            \spi_data_out_r_39__N_4511[22] , \spi_data_out_r_39__N_1404[22] , 
            \spi_data_out_r_39__N_1639[22] , \spi_data_out_r_39__N_1874[22] , 
            \spi_data_out_r_39__N_1169[22] , \spi_data_out_r_39__N_2109[22] , 
            \spi_data_out_r_39__N_934[22] , \spi_data_out_r_39__N_2344[22] , 
            \spi_data_out_r_39__N_5197[22] , \spi_data_out_r_39__N_4854[22] , 
            \spi_data_out_r[23] , \spi_data_out_r_39__N_3825[23] , \spi_data_out_r_39__N_4168[23] , 
            \spi_data_out_r_39__N_5540[23] , \spi_data_out_r_39__N_4511[23] , 
            \spi_data_out_r_39__N_1404[23] , \spi_data_out_r_39__N_1639[23] , 
            \spi_data_out_r_39__N_1874[23] , \spi_data_out_r_39__N_1169[23] , 
            \spi_data_out_r_39__N_2109[23] , \spi_data_out_r_39__N_934[23] , 
            \spi_data_out_r_39__N_2344[23] , \spi_data_out_r_39__N_5197[23] , 
            \spi_data_out_r_39__N_4854[23] , \spi_data_out_r[24] , \spi_data_out_r_39__N_3825[24] , 
            \spi_data_out_r_39__N_4168[24] , \spi_data_out_r_39__N_5540[24] , 
            \spi_data_out_r_39__N_4511[24] , \spi_data_out_r_39__N_1404[24] , 
            \spi_data_out_r_39__N_1639[24] , \spi_data_out_r_39__N_1874[24] , 
            \spi_data_out_r_39__N_1169[24] , \spi_data_out_r_39__N_2109[24] , 
            \spi_data_out_r_39__N_934[24] , \spi_data_out_r_39__N_2344[24] , 
            \spi_data_out_r_39__N_5197[24] , \spi_data_out_r_39__N_4854[24] , 
            \spi_data_out_r[25] , \spi_data_out_r_39__N_3825[25] , \spi_data_out_r_39__N_4168[25] , 
            \spi_data_out_r_39__N_5540[25] , \spi_data_out_r_39__N_4511[25] , 
            \spi_data_out_r_39__N_1404[25] , \spi_data_out_r_39__N_1639[25] , 
            \spi_data_out_r_39__N_1874[25] , \spi_data_out_r_39__N_1169[25] , 
            \spi_data_out_r_39__N_2109[25] , \spi_data_out_r_39__N_934[25] , 
            \spi_data_out_r_39__N_2344[25] , \spi_data_out_r_39__N_5197[25] , 
            \spi_data_out_r_39__N_4854[25] , \spi_data_out_r[26] , \spi_data_out_r_39__N_3825[26] , 
            \spi_data_out_r_39__N_4168[26] , \spi_data_out_r_39__N_5540[26] , 
            \spi_data_out_r_39__N_4511[26] , \spi_data_out_r_39__N_1404[26] , 
            \spi_data_out_r_39__N_1639[26] , \spi_data_out_r_39__N_1874[26] , 
            \spi_data_out_r_39__N_1169[26] , \spi_data_out_r_39__N_2109[26] , 
            \spi_data_out_r_39__N_934[26] , \spi_data_out_r_39__N_2344[26] , 
            \spi_data_out_r_39__N_5197[26] , \spi_data_out_r_39__N_4854[26] , 
            \spi_data_out_r[27] , \spi_data_out_r_39__N_3825[27] , \spi_data_out_r_39__N_4168[27] , 
            \spi_data_out_r_39__N_5540[27] , \spi_data_out_r_39__N_4511[27] , 
            \spi_data_out_r_39__N_1404[27] , \spi_data_out_r_39__N_1639[27] , 
            \spi_data_out_r_39__N_1874[27] , \spi_data_out_r_39__N_1169[27] , 
            \spi_data_out_r_39__N_2109[27] , \spi_data_out_r_39__N_934[27] , 
            \spi_data_out_r_39__N_2344[27] , \spi_data_out_r_39__N_5197[27] , 
            \spi_data_out_r_39__N_4854[27] , \spi_data_out_r[28] , \spi_data_out_r_39__N_3825[28] , 
            \spi_data_out_r_39__N_4168[28] , \spi_data_out_r_39__N_5540[28] , 
            \spi_data_out_r_39__N_4511[28] , \spi_data_out_r_39__N_1404[28] , 
            \spi_data_out_r_39__N_1639[28] , \spi_data_out_r_39__N_1874[28] , 
            \spi_data_out_r_39__N_1169[28] , \spi_data_out_r_39__N_2109[28] , 
            \spi_data_out_r_39__N_934[28] , \spi_data_out_r_39__N_2344[28] , 
            \spi_data_out_r_39__N_5197[28] , \spi_data_out_r_39__N_4854[28] , 
            \spi_data_out_r[29] , \spi_data_out_r_39__N_3825[29] , \spi_data_out_r_39__N_4168[29] , 
            \spi_data_out_r_39__N_5540[29] , \spi_data_out_r_39__N_4511[29] , 
            \spi_data_out_r_39__N_1404[29] , \spi_data_out_r_39__N_1639[29] , 
            \spi_data_out_r_39__N_1874[29] , \spi_data_out_r_39__N_1169[29] , 
            \spi_data_out_r_39__N_2109[29] , \spi_data_out_r_39__N_934[29] , 
            \spi_data_out_r_39__N_2344[29] , \spi_data_out_r_39__N_5197[29] , 
            \spi_data_out_r_39__N_4854[29] , n6, OW_ID_N_6182, \spi_data_out_r[30] , 
            \spi_data_out_r_39__N_3825[30] , \spi_data_out_r_39__N_4168[30] , 
            \spi_data_out_r_39__N_5540[30] , \spi_data_out_r_39__N_4511[30] , 
            \spi_data_out_r_39__N_1404[30] , \spi_data_out_r_39__N_1639[30] , 
            \spi_data_out_r_39__N_1874[30] , \spi_data_out_r_39__N_1169[30] , 
            \spi_data_out_r_39__N_2109[30] , \spi_data_out_r_39__N_934[30] , 
            \spi_data_out_r_39__N_2344[30] , \spi_data_out_r_39__N_5197[30] , 
            \spi_data_out_r_39__N_4854[30] , \spi_data_out_r[31] , \spi_data_out_r_39__N_3825[31] , 
            \spi_data_out_r_39__N_4168[31] , \spi_data_out_r_39__N_5540[31] , 
            \spi_data_out_r_39__N_4511[31] , \spi_data_out_r_39__N_1404[31] , 
            \spi_data_out_r_39__N_1639[31] , \spi_data_out_r_39__N_1874[31] , 
            \spi_data_out_r_39__N_1169[31] , \spi_data_out_r_39__N_2109[31] , 
            \spi_data_out_r_39__N_934[31] , \spi_data_out_r_39__N_2344[31] , 
            \spi_data_out_r_39__N_5197[31] , \spi_data_out_r_39__N_4854[31] , 
            \spi_data_out_r_39__N_4168[32] , \spi_data_out_r[32] , \spi_data_out_r_39__N_4854[32] , 
            \spi_data_out_r_39__N_5540[32] , \spi_data_out_r_39__N_4511[32] , 
            \spi_data_out_r_39__N_5197[32] , \spi_data_out_r_39__N_3825[32] , 
            \spi_data_out_r_39__N_4168[33] , \spi_data_out_r[33] , \spi_data_out_r_39__N_4854[33] , 
            \spi_data_out_r_39__N_5540[33] , \spi_data_out_r_39__N_4511[33] , 
            \spi_data_out_r_39__N_5197[33] , \spi_data_out_r_39__N_3825[33] , 
            \spi_data_out_r_39__N_4168[34] , \spi_data_out_r[34] , \spi_data_out_r_39__N_4854[34] , 
            \spi_data_out_r_39__N_5540[34] , \spi_data_out_r_39__N_4511[34] , 
            \spi_data_out_r_39__N_5197[34] , \spi_data_out_r_39__N_3825[34] , 
            \spi_data_out_r_39__N_4168[35] , \spi_data_out_r[35] , \spi_data_out_r_39__N_4854[35] , 
            \spi_data_out_r_39__N_5540[35] , \spi_data_out_r_39__N_4511[35] , 
            \spi_data_out_r_39__N_5197[35] , \spi_data_out_r_39__N_3825[35] , 
            \spi_data_out_r_39__N_4168[36] , \spi_data_out_r[36] , \spi_data_out_r_39__N_4854[36] , 
            \spi_data_out_r_39__N_5540[36] , \spi_data_out_r_39__N_4511[36] , 
            \spi_data_out_r_39__N_5197[36] , \spi_data_out_r_39__N_3825[36] , 
            \spi_data_out_r_39__N_4168[37] , \spi_data_out_r[37] , \spi_data_out_r_39__N_4854[37] , 
            \spi_data_out_r_39__N_5540[37] , \spi_data_out_r_39__N_4511[37] , 
            \spi_data_out_r_39__N_5197[37] , \spi_data_out_r_39__N_3825[37] , 
            \spi_data_out_r_39__N_4168[38] , \spi_data_out_r[38] , \spi_data_out_r_39__N_4854[38] , 
            \spi_data_out_r_39__N_5540[38] , \spi_data_out_r_39__N_4511[38] , 
            \spi_data_out_r_39__N_5197[38] , \spi_data_out_r_39__N_3825[38] , 
            \spi_data_out_r_39__N_4168[39] , \spi_data_out_r[39] , \spi_data_out_r_39__N_4854[39] , 
            \spi_data_out_r_39__N_5540[39] , \spi_data_out_r_39__N_4511[39] , 
            \spi_data_out_r_39__N_5197[39] , \spi_data_out_r_39__N_3825[39] , 
            \spi_data_out_r_39__N_5883[8] , \spi_data_out_r_39__N_5883[9] , 
            n47, \spi_data_out_r_39__N_3825[8] , n16, \spi_data_out_r_39__N_4511[8] , 
            n18, \spi_data_out_r_39__N_1639[8] , n5, \spi_data_out_r_39__N_1169[8] , 
            n3, \spi_data_out_r_39__N_3825[9] , n16_adj_1, \spi_data_out_r_39__N_5540[9] , 
            n21, \spi_data_out_r_39__N_1639[9] , n5_adj_2, \spi_data_out_r_39__N_934[9] , 
            n2, n30165, \spi_data_out_r_39__N_5540[2] , n21_adj_3, \spi_data_out_r_39__N_4854[2] , 
            n19, GND_net, \spi_data_out_r_39__N_2109[2] , n7, n22, 
            \spi_data_out_r_39__N_2934[2] , clear_intrpt, n14, \spi_data_out_r_39__N_2579[2] , 
            clear_intrpt_adj_4, n9, \spi_data_out_r[0] , \spi_data_out_r_39__N_4854[0] , 
            \spi_data_out_r_39__N_4168[0] , \spi_data_out_r_39__N_5197[0] , 
            \spi_data_out_r_39__N_2650[0] , clear_intrpt_adj_5, \spi_data_out_r_39__N_2863[0] , 
            clear_intrpt_adj_6, \spi_data_out_r_39__N_2934[0] , \spi_data_out_r_39__N_770[0] , 
            spi_data_out_r_39__N_810, \spi_data_out_r_39__N_3005[0] , clear_intrpt_adj_7, 
            \spi_data_out_r_39__N_2109[0] , \spi_data_out_r_39__N_3825[0] , 
            \spi_data_out_r_39__N_5540[0] , \spi_data_out_r_39__N_2344[0] , 
            \spi_data_out_r_39__N_934[0] , \spi_data_out_r_39__N_1404[0] , 
            \spi_data_out_r_39__N_1639[0] , \spi_data_out_r_39__N_1169[0] , 
            \spi_data_out_r_39__N_1874[0] , \spi_data_out_r_39__N_4511[0] , 
            \spi_data_out_r_39__N_2792[0] , \spi_data_out_r_39__N_2579[0] , 
            clear_intrpt_adj_8, \spi_data_out_r_39__N_2721[0] , clear_intrpt_adj_9, 
            \uart_slot_en[3] , pin_io_out_65, n24700, pin_io_c_68, \quad_a[6] , 
            pin_io_out_69, \quad_b[6] , UC_TXD0_c, OW_ID_N_6176, n30083, 
            pin_io_c_63, \pin_intrpt[19] , pin_io_c_64, \pin_intrpt[20] , 
            pin_io_c_62, \pin_intrpt[18] , n7258, \quad_homing[0] , 
            n25889, \spi_data_out_r[1] , \spi_data_out_r_39__N_2934[1] , 
            \spi_data_out_r_39__N_4511[1] , \spi_data_out_r_39__N_5197[1] , 
            \spi_data_out_r_39__N_3825[1] , \spi_data_out_r_39__N_2863[1] , 
            \spi_data_out_r_39__N_3005[1] , \spi_data_out_r_39__N_2579[1] , 
            \spi_data_out_r_39__N_2792[1] , \spi_data_out_r_39__N_2650[1] , 
            \spi_data_out_r_39__N_2721[1] , \spi_data_out_r_39__N_1169[1] , 
            \spi_data_out_r_39__N_4168[1] , \spi_data_out_r_39__N_5540[1] , 
            \spi_data_out_r_39__N_2344[1] , \spi_data_out_r_39__N_1639[1] , 
            \spi_data_out_r_39__N_934[1] , \spi_data_out_r_39__N_2109[1] , 
            \spi_data_out_r_39__N_1404[1] , \spi_data_out_r_39__N_1874[1] , 
            \spi_data_out_r_39__N_4854[1] , \spi_data_out_r[3] , \spi_data_out_r_39__N_3825[3] , 
            \spi_data_out_r_39__N_4168[3] , \spi_data_out_r_39__N_5540[3] , 
            \spi_data_out_r_39__N_4511[3] , \spi_data_out_r_39__N_1404[3] , 
            \spi_data_out_r_39__N_1639[3] , \spi_data_out_r_39__N_1874[3] , 
            \spi_data_out_r_39__N_1169[3] , \spi_data_out_r_39__N_2109[3] , 
            \spi_data_out_r_39__N_934[3] , \spi_data_out_r_39__N_2344[3] , 
            \spi_data_out_r_39__N_5197[3] , \spi_data_out_r_39__N_4854[3] , 
            \spi_data_out_r[4] , \spi_data_out_r_39__N_3825[4] , \spi_data_out_r_39__N_4168[4] , 
            ENC_O_N_6184) /* synthesis syn_module_defined=1 */ ;
    input \spi_data_out_r_39__N_5540[4] ;
    input spi_data_out_r_39__N_5580;
    input \spi_data_out_r_39__N_4511[4] ;
    input spi_data_out_r_39__N_4551;
    input clk;
    input \spi_data_out_r_39__N_1404[4] ;
    input \spi_data_out_r_39__N_1639[4] ;
    input spi_data_out_r_39__N_1444;
    input spi_data_out_r_39__N_1679;
    input \spi_data_out_r_39__N_1874[4] ;
    input spi_data_out_r_39__N_1914;
    input \spi_data_out_r_39__N_1169[4] ;
    input spi_data_out_r_39__N_1209;
    input \spi_data_out_r_39__N_2109[4] ;
    input \spi_data_out_r_39__N_934[4] ;
    input spi_data_out_r_39__N_2149;
    input spi_data_out_r_39__N_974;
    input \spi_data_out_r_39__N_2344[4] ;
    input spi_data_out_r_39__N_2384;
    input \spi_data_out_r_39__N_5197[4] ;
    input \spi_data_out_r_39__N_4854[4] ;
    input spi_data_out_r_39__N_5237;
    input spi_data_out_r_39__N_4894;
    output spi_data_out_r_39__N_5923;
    output \spi_data_out_r[5] ;
    input \spi_data_out_r_39__N_3825[5] ;
    input \spi_data_out_r_39__N_4168[5] ;
    input spi_data_out_r_39__N_3865;
    input spi_data_out_r_39__N_4208;
    input \spi_data_out_r_39__N_5540[5] ;
    output reset_r;
    input n30185;
    input n30028;
    output NSL;
    input clk_1MHz;
    input \spi_data_out_r_39__N_4511[5] ;
    input \spi_data_out_r_39__N_1404[5] ;
    input \spi_data_out_r_39__N_1639[5] ;
    input \spi_data_out_r_39__N_1874[5] ;
    input \spi_data_out_r_39__N_1169[5] ;
    input \spi_data_out_r_39__N_2109[5] ;
    input \spi_data_out_r_39__N_934[5] ;
    input \spi_data_out_r_39__N_2344[5] ;
    input \spi_data_out_r_39__N_5197[5] ;
    input \spi_data_out_r_39__N_4854[5] ;
    input clk_enable_180;
    input \spi_data_r[0] ;
    output \spi_data_out_r[6] ;
    input \spi_data_out_r_39__N_3825[6] ;
    input \spi_data_out_r_39__N_4168[6] ;
    input \spi_data_out_r_39__N_5540[6] ;
    input \spi_data_out_r_39__N_4511[6] ;
    input \spi_data_out_r_39__N_1404[6] ;
    input \spi_data_out_r_39__N_1639[6] ;
    input \spi_data_out_r_39__N_1874[6] ;
    input \spi_data_out_r_39__N_1169[6] ;
    input \spi_data_out_r_39__N_2109[6] ;
    input \spi_data_out_r_39__N_934[6] ;
    input \spi_data_out_r_39__N_2344[6] ;
    input \spi_data_out_r_39__N_5197[6] ;
    input \spi_data_out_r_39__N_4854[6] ;
    output \spi_data_out_r[7] ;
    input \spi_data_out_r_39__N_3825[7] ;
    input \spi_data_out_r_39__N_4168[7] ;
    input \spi_data_out_r_39__N_5540[7] ;
    input \spi_data_out_r_39__N_4511[7] ;
    input \spi_data_out_r_39__N_1404[7] ;
    input \spi_data_out_r_39__N_1639[7] ;
    output n30143;
    input \spi_data_out_r_39__N_1874[7] ;
    input \spi_data_out_r_39__N_1169[7] ;
    input \spi_data_out_r_39__N_2109[7] ;
    input \spi_data_out_r_39__N_934[7] ;
    input \spi_data_out_r_39__N_2344[7] ;
    input \spi_data_out_r_39__N_5197[7] ;
    input \spi_data_out_r_39__N_4854[7] ;
    input resetn_c;
    output \spi_data_out_r[10] ;
    input \spi_data_out_r_39__N_3825[10] ;
    input \spi_data_out_r_39__N_4168[10] ;
    input \spi_data_r[2] ;
    input \spi_data_r[1] ;
    input \spi_data_out_r_39__N_5540[10] ;
    input \spi_data_out_r_39__N_4511[10] ;
    input \spi_data_out_r_39__N_1404[10] ;
    input \spi_data_out_r_39__N_1639[10] ;
    input \spi_data_out_r_39__N_1874[10] ;
    input \spi_data_out_r_39__N_1169[10] ;
    input \spi_data_out_r_39__N_2109[10] ;
    input \spi_data_out_r_39__N_934[10] ;
    input \spi_data_out_r_39__N_2344[10] ;
    input \spi_data_out_r_39__N_5197[10] ;
    input \spi_data_out_r_39__N_4854[10] ;
    output \spi_data_out_r[11] ;
    input \spi_data_out_r_39__N_3825[11] ;
    input \spi_data_out_r_39__N_4168[11] ;
    input \spi_data_out_r_39__N_5540[11] ;
    input \spi_data_out_r_39__N_4511[11] ;
    input \spi_data_out_r_39__N_1404[11] ;
    input \spi_data_out_r_39__N_1639[11] ;
    input \spi_data_out_r_39__N_1874[11] ;
    input \spi_data_out_r_39__N_1169[11] ;
    input \spi_data_out_r_39__N_2109[11] ;
    input \spi_data_out_r_39__N_934[11] ;
    input \spi_data_out_r_39__N_2344[11] ;
    input \spi_data_out_r_39__N_5197[11] ;
    input \spi_data_out_r_39__N_4854[11] ;
    output \spi_data_out_r[12] ;
    input \spi_data_out_r_39__N_3825[12] ;
    input \spi_data_out_r_39__N_4168[12] ;
    input \spi_data_out_r_39__N_5540[12] ;
    input \spi_data_out_r_39__N_4511[12] ;
    input \spi_data_out_r_39__N_1404[12] ;
    input \spi_data_out_r_39__N_1639[12] ;
    input \spi_data_out_r_39__N_1874[12] ;
    input \spi_data_out_r_39__N_1169[12] ;
    input \spi_data_out_r_39__N_2109[12] ;
    input \spi_data_out_r_39__N_934[12] ;
    input \spi_data_out_r_39__N_2344[12] ;
    input \spi_data_out_r_39__N_5197[12] ;
    input \spi_data_out_r_39__N_4854[12] ;
    output \spi_data_out_r[13] ;
    input \spi_data_out_r_39__N_3825[13] ;
    input \spi_data_out_r_39__N_4168[13] ;
    output digital_output_r;
    input clk_enable_222;
    input n28550;
    input \spi_data_out_r_39__N_5540[13] ;
    input EM_STOP;
    input n25741;
    input n23916;
    input \spi_data_out_r_39__N_4511[13] ;
    input \spi_data_out_r_39__N_1404[13] ;
    input \spi_data_out_r_39__N_1639[13] ;
    input \spi_data_out_r_39__N_1874[13] ;
    input \spi_data_out_r_39__N_1169[13] ;
    input \spi_data_out_r_39__N_2109[13] ;
    input \spi_data_out_r_39__N_934[13] ;
    input \spi_data_out_r_39__N_2344[13] ;
    input \spi_data_out_r_39__N_5197[13] ;
    input \spi_data_out_r_39__N_4854[13] ;
    output \spi_data_out_r[14] ;
    input \spi_data_out_r_39__N_3825[14] ;
    input \spi_data_out_r_39__N_4168[14] ;
    input \spi_data_out_r_39__N_5540[14] ;
    input \spi_data_out_r_39__N_4511[14] ;
    input \spi_data_out_r_39__N_1404[14] ;
    input \spi_data_out_r_39__N_1639[14] ;
    input \spi_data_out_r_39__N_1874[14] ;
    input \spi_data_out_r_39__N_1169[14] ;
    input \spi_data_out_r_39__N_2109[14] ;
    input \spi_data_out_r_39__N_934[14] ;
    input \spi_data_out_r_39__N_2344[14] ;
    input \spi_data_out_r_39__N_5197[14] ;
    input \spi_data_out_r_39__N_4854[14] ;
    output \spi_data_out_r[15] ;
    input \spi_data_out_r_39__N_3825[15] ;
    input \spi_data_out_r_39__N_4168[15] ;
    input \spi_data_out_r_39__N_5540[15] ;
    input \spi_data_out_r_39__N_4511[15] ;
    input \spi_data_out_r_39__N_1404[15] ;
    input \spi_data_out_r_39__N_1639[15] ;
    input \spi_data_out_r_39__N_1874[15] ;
    input \spi_data_out_r_39__N_1169[15] ;
    input \spi_data_out_r_39__N_2109[15] ;
    input \spi_data_out_r_39__N_934[15] ;
    input \spi_data_out_r_39__N_2344[15] ;
    input \spi_data_out_r_39__N_5197[15] ;
    input \spi_data_out_r_39__N_4854[15] ;
    output \spi_data_out_r[16] ;
    input \spi_data_out_r_39__N_3825[16] ;
    input \spi_data_out_r_39__N_4168[16] ;
    input \spi_data_out_r_39__N_5540[16] ;
    input \spi_data_out_r_39__N_4511[16] ;
    input \spi_data_out_r_39__N_1404[16] ;
    input \spi_data_out_r_39__N_1639[16] ;
    input \spi_data_out_r_39__N_1874[16] ;
    input \spi_data_out_r_39__N_1169[16] ;
    input \spi_data_out_r_39__N_2109[16] ;
    input \spi_data_out_r_39__N_934[16] ;
    input \spi_data_out_r_39__N_2344[16] ;
    input \spi_data_out_r_39__N_5197[16] ;
    input \spi_data_out_r_39__N_4854[16] ;
    output \spi_data_out_r[17] ;
    input \spi_data_out_r_39__N_3825[17] ;
    input \spi_data_out_r_39__N_4168[17] ;
    input \spi_data_out_r_39__N_5540[17] ;
    input \spi_data_out_r_39__N_4511[17] ;
    input \spi_data_out_r_39__N_1404[17] ;
    input \spi_data_out_r_39__N_1639[17] ;
    input spi_data_out_r_39__N_6220;
    input \spi_data_out_r_39__N_1874[17] ;
    input \spi_data_out_r_39__N_1169[17] ;
    input \spi_data_out_r_39__N_2109[17] ;
    input \spi_data_out_r_39__N_934[17] ;
    input \spi_data_out_r_39__N_2344[17] ;
    input \spi_data_out_r_39__N_5197[17] ;
    input \spi_data_out_r_39__N_4854[17] ;
    output \spi_data_out_r[18] ;
    input \spi_data_out_r_39__N_3825[18] ;
    input \spi_data_out_r_39__N_4168[18] ;
    input \spi_data_out_r_39__N_5540[18] ;
    input \spi_data_out_r_39__N_4511[18] ;
    input \spi_data_out_r_39__N_1404[18] ;
    input \spi_data_out_r_39__N_1639[18] ;
    input \spi_data_out_r_39__N_1874[18] ;
    input \spi_data_out_r_39__N_1169[18] ;
    input \spi_data_out_r_39__N_2109[18] ;
    input \spi_data_out_r_39__N_934[18] ;
    input \spi_data_out_r_39__N_2344[18] ;
    input \spi_data_out_r_39__N_5197[18] ;
    input \spi_data_out_r_39__N_4854[18] ;
    output \spi_data_out_r[19] ;
    input \spi_data_out_r_39__N_3825[19] ;
    input \spi_data_out_r_39__N_4168[19] ;
    input \spi_data_out_r_39__N_5540[19] ;
    input \spi_data_out_r_39__N_4511[19] ;
    input \spi_data_out_r_39__N_1404[19] ;
    input \spi_data_out_r_39__N_1639[19] ;
    input \spi_data_out_r_39__N_1874[19] ;
    input \spi_data_out_r_39__N_1169[19] ;
    input \spi_data_out_r_39__N_2109[19] ;
    input \spi_data_out_r_39__N_934[19] ;
    input \spi_data_out_r_39__N_2344[19] ;
    input \spi_data_out_r_39__N_5197[19] ;
    input \spi_data_out_r_39__N_4854[19] ;
    output \spi_data_out_r[20] ;
    input \spi_data_out_r_39__N_3825[20] ;
    input \spi_data_out_r_39__N_4168[20] ;
    input \spi_data_out_r_39__N_5540[20] ;
    input \spi_data_out_r_39__N_4511[20] ;
    input \spi_data_out_r_39__N_1404[20] ;
    input \spi_data_out_r_39__N_1639[20] ;
    input \spi_data_out_r_39__N_1874[20] ;
    input \spi_data_out_r_39__N_1169[20] ;
    input \spi_data_out_r_39__N_2109[20] ;
    input \spi_data_out_r_39__N_934[20] ;
    input \spi_data_out_r_39__N_2344[20] ;
    input \spi_data_out_r_39__N_5197[20] ;
    input \spi_data_out_r_39__N_4854[20] ;
    output \spi_data_out_r[21] ;
    input \spi_data_out_r_39__N_3825[21] ;
    input \spi_data_out_r_39__N_4168[21] ;
    input \spi_data_out_r_39__N_5540[21] ;
    input \spi_data_out_r_39__N_4511[21] ;
    input \spi_data_out_r_39__N_1404[21] ;
    input \spi_data_out_r_39__N_1639[21] ;
    input \spi_data_out_r_39__N_1874[21] ;
    input \spi_data_out_r_39__N_1169[21] ;
    input \spi_data_out_r_39__N_2109[21] ;
    input \spi_data_out_r_39__N_934[21] ;
    input \spi_data_out_r_39__N_2344[21] ;
    input \spi_data_out_r_39__N_5197[21] ;
    input \spi_data_out_r_39__N_4854[21] ;
    output \spi_data_out_r[22] ;
    input \spi_data_out_r_39__N_3825[22] ;
    input \spi_data_out_r_39__N_4168[22] ;
    input \spi_data_out_r_39__N_5540[22] ;
    input \spi_data_out_r_39__N_4511[22] ;
    input \spi_data_out_r_39__N_1404[22] ;
    input \spi_data_out_r_39__N_1639[22] ;
    input \spi_data_out_r_39__N_1874[22] ;
    input \spi_data_out_r_39__N_1169[22] ;
    input \spi_data_out_r_39__N_2109[22] ;
    input \spi_data_out_r_39__N_934[22] ;
    input \spi_data_out_r_39__N_2344[22] ;
    input \spi_data_out_r_39__N_5197[22] ;
    input \spi_data_out_r_39__N_4854[22] ;
    output \spi_data_out_r[23] ;
    input \spi_data_out_r_39__N_3825[23] ;
    input \spi_data_out_r_39__N_4168[23] ;
    input \spi_data_out_r_39__N_5540[23] ;
    input \spi_data_out_r_39__N_4511[23] ;
    input \spi_data_out_r_39__N_1404[23] ;
    input \spi_data_out_r_39__N_1639[23] ;
    input \spi_data_out_r_39__N_1874[23] ;
    input \spi_data_out_r_39__N_1169[23] ;
    input \spi_data_out_r_39__N_2109[23] ;
    input \spi_data_out_r_39__N_934[23] ;
    input \spi_data_out_r_39__N_2344[23] ;
    input \spi_data_out_r_39__N_5197[23] ;
    input \spi_data_out_r_39__N_4854[23] ;
    output \spi_data_out_r[24] ;
    input \spi_data_out_r_39__N_3825[24] ;
    input \spi_data_out_r_39__N_4168[24] ;
    input \spi_data_out_r_39__N_5540[24] ;
    input \spi_data_out_r_39__N_4511[24] ;
    input \spi_data_out_r_39__N_1404[24] ;
    input \spi_data_out_r_39__N_1639[24] ;
    input \spi_data_out_r_39__N_1874[24] ;
    input \spi_data_out_r_39__N_1169[24] ;
    input \spi_data_out_r_39__N_2109[24] ;
    input \spi_data_out_r_39__N_934[24] ;
    input \spi_data_out_r_39__N_2344[24] ;
    input \spi_data_out_r_39__N_5197[24] ;
    input \spi_data_out_r_39__N_4854[24] ;
    output \spi_data_out_r[25] ;
    input \spi_data_out_r_39__N_3825[25] ;
    input \spi_data_out_r_39__N_4168[25] ;
    input \spi_data_out_r_39__N_5540[25] ;
    input \spi_data_out_r_39__N_4511[25] ;
    input \spi_data_out_r_39__N_1404[25] ;
    input \spi_data_out_r_39__N_1639[25] ;
    input \spi_data_out_r_39__N_1874[25] ;
    input \spi_data_out_r_39__N_1169[25] ;
    input \spi_data_out_r_39__N_2109[25] ;
    input \spi_data_out_r_39__N_934[25] ;
    input \spi_data_out_r_39__N_2344[25] ;
    input \spi_data_out_r_39__N_5197[25] ;
    input \spi_data_out_r_39__N_4854[25] ;
    output \spi_data_out_r[26] ;
    input \spi_data_out_r_39__N_3825[26] ;
    input \spi_data_out_r_39__N_4168[26] ;
    input \spi_data_out_r_39__N_5540[26] ;
    input \spi_data_out_r_39__N_4511[26] ;
    input \spi_data_out_r_39__N_1404[26] ;
    input \spi_data_out_r_39__N_1639[26] ;
    input \spi_data_out_r_39__N_1874[26] ;
    input \spi_data_out_r_39__N_1169[26] ;
    input \spi_data_out_r_39__N_2109[26] ;
    input \spi_data_out_r_39__N_934[26] ;
    input \spi_data_out_r_39__N_2344[26] ;
    input \spi_data_out_r_39__N_5197[26] ;
    input \spi_data_out_r_39__N_4854[26] ;
    output \spi_data_out_r[27] ;
    input \spi_data_out_r_39__N_3825[27] ;
    input \spi_data_out_r_39__N_4168[27] ;
    input \spi_data_out_r_39__N_5540[27] ;
    input \spi_data_out_r_39__N_4511[27] ;
    input \spi_data_out_r_39__N_1404[27] ;
    input \spi_data_out_r_39__N_1639[27] ;
    input \spi_data_out_r_39__N_1874[27] ;
    input \spi_data_out_r_39__N_1169[27] ;
    input \spi_data_out_r_39__N_2109[27] ;
    input \spi_data_out_r_39__N_934[27] ;
    input \spi_data_out_r_39__N_2344[27] ;
    input \spi_data_out_r_39__N_5197[27] ;
    input \spi_data_out_r_39__N_4854[27] ;
    output \spi_data_out_r[28] ;
    input \spi_data_out_r_39__N_3825[28] ;
    input \spi_data_out_r_39__N_4168[28] ;
    input \spi_data_out_r_39__N_5540[28] ;
    input \spi_data_out_r_39__N_4511[28] ;
    input \spi_data_out_r_39__N_1404[28] ;
    input \spi_data_out_r_39__N_1639[28] ;
    input \spi_data_out_r_39__N_1874[28] ;
    input \spi_data_out_r_39__N_1169[28] ;
    input \spi_data_out_r_39__N_2109[28] ;
    input \spi_data_out_r_39__N_934[28] ;
    input \spi_data_out_r_39__N_2344[28] ;
    input \spi_data_out_r_39__N_5197[28] ;
    input \spi_data_out_r_39__N_4854[28] ;
    output \spi_data_out_r[29] ;
    input \spi_data_out_r_39__N_3825[29] ;
    input \spi_data_out_r_39__N_4168[29] ;
    input \spi_data_out_r_39__N_5540[29] ;
    input \spi_data_out_r_39__N_4511[29] ;
    input \spi_data_out_r_39__N_1404[29] ;
    input \spi_data_out_r_39__N_1639[29] ;
    input \spi_data_out_r_39__N_1874[29] ;
    input \spi_data_out_r_39__N_1169[29] ;
    input \spi_data_out_r_39__N_2109[29] ;
    input \spi_data_out_r_39__N_934[29] ;
    input \spi_data_out_r_39__N_2344[29] ;
    input \spi_data_out_r_39__N_5197[29] ;
    input \spi_data_out_r_39__N_4854[29] ;
    input n6;
    output OW_ID_N_6182;
    output \spi_data_out_r[30] ;
    input \spi_data_out_r_39__N_3825[30] ;
    input \spi_data_out_r_39__N_4168[30] ;
    input \spi_data_out_r_39__N_5540[30] ;
    input \spi_data_out_r_39__N_4511[30] ;
    input \spi_data_out_r_39__N_1404[30] ;
    input \spi_data_out_r_39__N_1639[30] ;
    input \spi_data_out_r_39__N_1874[30] ;
    input \spi_data_out_r_39__N_1169[30] ;
    input \spi_data_out_r_39__N_2109[30] ;
    input \spi_data_out_r_39__N_934[30] ;
    input \spi_data_out_r_39__N_2344[30] ;
    input \spi_data_out_r_39__N_5197[30] ;
    input \spi_data_out_r_39__N_4854[30] ;
    output \spi_data_out_r[31] ;
    input \spi_data_out_r_39__N_3825[31] ;
    input \spi_data_out_r_39__N_4168[31] ;
    input \spi_data_out_r_39__N_5540[31] ;
    input \spi_data_out_r_39__N_4511[31] ;
    input \spi_data_out_r_39__N_1404[31] ;
    input \spi_data_out_r_39__N_1639[31] ;
    input \spi_data_out_r_39__N_1874[31] ;
    input \spi_data_out_r_39__N_1169[31] ;
    input \spi_data_out_r_39__N_2109[31] ;
    input \spi_data_out_r_39__N_934[31] ;
    input \spi_data_out_r_39__N_2344[31] ;
    input \spi_data_out_r_39__N_5197[31] ;
    input \spi_data_out_r_39__N_4854[31] ;
    input \spi_data_out_r_39__N_4168[32] ;
    output \spi_data_out_r[32] ;
    input \spi_data_out_r_39__N_4854[32] ;
    input \spi_data_out_r_39__N_5540[32] ;
    input \spi_data_out_r_39__N_4511[32] ;
    input \spi_data_out_r_39__N_5197[32] ;
    input \spi_data_out_r_39__N_3825[32] ;
    input \spi_data_out_r_39__N_4168[33] ;
    output \spi_data_out_r[33] ;
    input \spi_data_out_r_39__N_4854[33] ;
    input \spi_data_out_r_39__N_5540[33] ;
    input \spi_data_out_r_39__N_4511[33] ;
    input \spi_data_out_r_39__N_5197[33] ;
    input \spi_data_out_r_39__N_3825[33] ;
    input \spi_data_out_r_39__N_4168[34] ;
    output \spi_data_out_r[34] ;
    input \spi_data_out_r_39__N_4854[34] ;
    input \spi_data_out_r_39__N_5540[34] ;
    input \spi_data_out_r_39__N_4511[34] ;
    input \spi_data_out_r_39__N_5197[34] ;
    input \spi_data_out_r_39__N_3825[34] ;
    input \spi_data_out_r_39__N_4168[35] ;
    output \spi_data_out_r[35] ;
    input \spi_data_out_r_39__N_4854[35] ;
    input \spi_data_out_r_39__N_5540[35] ;
    input \spi_data_out_r_39__N_4511[35] ;
    input \spi_data_out_r_39__N_5197[35] ;
    input \spi_data_out_r_39__N_3825[35] ;
    input \spi_data_out_r_39__N_4168[36] ;
    output \spi_data_out_r[36] ;
    input \spi_data_out_r_39__N_4854[36] ;
    input \spi_data_out_r_39__N_5540[36] ;
    input \spi_data_out_r_39__N_4511[36] ;
    input \spi_data_out_r_39__N_5197[36] ;
    input \spi_data_out_r_39__N_3825[36] ;
    input \spi_data_out_r_39__N_4168[37] ;
    output \spi_data_out_r[37] ;
    input \spi_data_out_r_39__N_4854[37] ;
    input \spi_data_out_r_39__N_5540[37] ;
    input \spi_data_out_r_39__N_4511[37] ;
    input \spi_data_out_r_39__N_5197[37] ;
    input \spi_data_out_r_39__N_3825[37] ;
    input \spi_data_out_r_39__N_4168[38] ;
    output \spi_data_out_r[38] ;
    input \spi_data_out_r_39__N_4854[38] ;
    input \spi_data_out_r_39__N_5540[38] ;
    input \spi_data_out_r_39__N_4511[38] ;
    input \spi_data_out_r_39__N_5197[38] ;
    input \spi_data_out_r_39__N_3825[38] ;
    input \spi_data_out_r_39__N_4168[39] ;
    output \spi_data_out_r[39] ;
    input \spi_data_out_r_39__N_4854[39] ;
    input \spi_data_out_r_39__N_5540[39] ;
    input \spi_data_out_r_39__N_4511[39] ;
    input \spi_data_out_r_39__N_5197[39] ;
    input \spi_data_out_r_39__N_3825[39] ;
    output \spi_data_out_r_39__N_5883[8] ;
    output \spi_data_out_r_39__N_5883[9] ;
    input n47;
    input \spi_data_out_r_39__N_3825[8] ;
    output n16;
    input \spi_data_out_r_39__N_4511[8] ;
    output n18;
    input \spi_data_out_r_39__N_1639[8] ;
    output n5;
    input \spi_data_out_r_39__N_1169[8] ;
    output n3;
    input \spi_data_out_r_39__N_3825[9] ;
    output n16_adj_1;
    input \spi_data_out_r_39__N_5540[9] ;
    output n21;
    input \spi_data_out_r_39__N_1639[9] ;
    output n5_adj_2;
    input \spi_data_out_r_39__N_934[9] ;
    output n2;
    output n30165;
    input \spi_data_out_r_39__N_5540[2] ;
    output n21_adj_3;
    input \spi_data_out_r_39__N_4854[2] ;
    output n19;
    input GND_net;
    input \spi_data_out_r_39__N_2109[2] ;
    output n7;
    output n22;
    input \spi_data_out_r_39__N_2934[2] ;
    input clear_intrpt;
    output n14;
    input \spi_data_out_r_39__N_2579[2] ;
    input clear_intrpt_adj_4;
    output n9;
    output \spi_data_out_r[0] ;
    input \spi_data_out_r_39__N_4854[0] ;
    input \spi_data_out_r_39__N_4168[0] ;
    input \spi_data_out_r_39__N_5197[0] ;
    input \spi_data_out_r_39__N_2650[0] ;
    input clear_intrpt_adj_5;
    input \spi_data_out_r_39__N_2863[0] ;
    input clear_intrpt_adj_6;
    input \spi_data_out_r_39__N_2934[0] ;
    input \spi_data_out_r_39__N_770[0] ;
    input spi_data_out_r_39__N_810;
    input \spi_data_out_r_39__N_3005[0] ;
    input clear_intrpt_adj_7;
    input \spi_data_out_r_39__N_2109[0] ;
    input \spi_data_out_r_39__N_3825[0] ;
    input \spi_data_out_r_39__N_5540[0] ;
    input \spi_data_out_r_39__N_2344[0] ;
    input \spi_data_out_r_39__N_934[0] ;
    input \spi_data_out_r_39__N_1404[0] ;
    input \spi_data_out_r_39__N_1639[0] ;
    input \spi_data_out_r_39__N_1169[0] ;
    input \spi_data_out_r_39__N_1874[0] ;
    input \spi_data_out_r_39__N_4511[0] ;
    input \spi_data_out_r_39__N_2792[0] ;
    input \spi_data_out_r_39__N_2579[0] ;
    input clear_intrpt_adj_8;
    input \spi_data_out_r_39__N_2721[0] ;
    input clear_intrpt_adj_9;
    input \uart_slot_en[3] ;
    input pin_io_out_65;
    output n24700;
    input pin_io_c_68;
    output \quad_a[6] ;
    input pin_io_out_69;
    output \quad_b[6] ;
    input UC_TXD0_c;
    output OW_ID_N_6176;
    output n30083;
    input pin_io_c_63;
    output \pin_intrpt[19] ;
    input pin_io_c_64;
    output \pin_intrpt[20] ;
    input pin_io_c_62;
    output \pin_intrpt[18] ;
    output n7258;
    input \quad_homing[0] ;
    output n25889;
    output \spi_data_out_r[1] ;
    input \spi_data_out_r_39__N_2934[1] ;
    input \spi_data_out_r_39__N_4511[1] ;
    input \spi_data_out_r_39__N_5197[1] ;
    input \spi_data_out_r_39__N_3825[1] ;
    input \spi_data_out_r_39__N_2863[1] ;
    input \spi_data_out_r_39__N_3005[1] ;
    input \spi_data_out_r_39__N_2579[1] ;
    input \spi_data_out_r_39__N_2792[1] ;
    input \spi_data_out_r_39__N_2650[1] ;
    input \spi_data_out_r_39__N_2721[1] ;
    input \spi_data_out_r_39__N_1169[1] ;
    input \spi_data_out_r_39__N_4168[1] ;
    input \spi_data_out_r_39__N_5540[1] ;
    input \spi_data_out_r_39__N_2344[1] ;
    input \spi_data_out_r_39__N_1639[1] ;
    input \spi_data_out_r_39__N_934[1] ;
    input \spi_data_out_r_39__N_2109[1] ;
    input \spi_data_out_r_39__N_1404[1] ;
    input \spi_data_out_r_39__N_1874[1] ;
    input \spi_data_out_r_39__N_4854[1] ;
    output \spi_data_out_r[3] ;
    input \spi_data_out_r_39__N_3825[3] ;
    input \spi_data_out_r_39__N_4168[3] ;
    input \spi_data_out_r_39__N_5540[3] ;
    input \spi_data_out_r_39__N_4511[3] ;
    input \spi_data_out_r_39__N_1404[3] ;
    input \spi_data_out_r_39__N_1639[3] ;
    input \spi_data_out_r_39__N_1874[3] ;
    input \spi_data_out_r_39__N_1169[3] ;
    input \spi_data_out_r_39__N_2109[3] ;
    input \spi_data_out_r_39__N_934[3] ;
    input \spi_data_out_r_39__N_2344[3] ;
    input \spi_data_out_r_39__N_5197[3] ;
    input \spi_data_out_r_39__N_4854[3] ;
    output \spi_data_out_r[4] ;
    input \spi_data_out_r_39__N_3825[4] ;
    input \spi_data_out_r_39__N_4168[4] ;
    output ENC_O_N_6184;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    wire clk_1MHz /* synthesis SET_AS_NETWORK=clk_1MHz, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(136[6:14])
    wire \pin_intrpt[20]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[20] */ ;   // c:/s_links/sources/mcm_top.v(93[46:56])
    
    wire n27971, n3_c, n27977, n27967, n22_c, n27975;
    wire [51:0]SLO_buf;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire SLO_buf_51__N_6073;
    wire [51:0]SLO;   // c:/s_links/sources/slot_cards/stepper.v(63[12:15])
    
    wire n27961, n27957, n8;
    wire [39:0]spi_data_out_r_39__N_5883;
    
    wire n27681, n27689, n27687, n27673, n27683, n3_adj_6595, clk_enable_46, 
        clk_1MHz_enable_9, NSL_N_6215, n27679, n22_adj_6596, n27669, 
        n8_adj_6597;
    wire [2:0]mode;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    wire n28065, n28073, n28071, n28057, n28067, n3_adj_6598, n28063, 
        n22_adj_6599, n28053, n8_adj_6600, prev_MA_Temp, MA_Temp, 
        n27729, n27737, n27735, n27721, n27731, n3_adj_6601, n27727, 
        n22_adj_6602, prev_MA;
    wire [39:0]spi_data_out_r_39__N_6134;
    wire [7:0]Cnt;   // c:/s_links/sources/slot_cards/stepper.v(62[11:14])
    
    wire clk_1MHz_enable_49;
    wire [7:0]n199;
    
    wire n27717, n8_adj_6603;
    wire [11:0]n93;
    wire [11:0]n53;
    
    wire n27585, n27593, n27591, n27577, n27587, n3_adj_6604, n27583, 
        n22_adj_6605, n27573, n8_adj_6606, n27849, n27857, n27855, 
        n27841, n27851, n3_adj_6607, n27847, n22_adj_6608, n27837, 
        n8_adj_6609, n28089, n28097, n28095, n28081, n28091, n3_adj_6610, 
        n28087, n22_adj_6611, n28077, n8_adj_6612, n27561, n27569, 
        n27567, n27553, n27563, n3_adj_6613, n27559, n22_adj_6614, 
        n27549, n8_adj_6615, n28041, n28049, n28047, n28033, n28043, 
        n3_adj_6616, n28039, n22_adj_6617, n28029, n8_adj_6618, n27801, 
        n27809, n27807, n27793, n27803, n3_adj_6619, n27799, n22_adj_6620, 
        n27789, n8_adj_6621, n28017, n28025, n28023, n28009, n28019, 
        n3_adj_6622, n18534, n30164, n29680, n28015, n22_adj_6623, 
        n28005, n8_adj_6624, n28113, n28121, n28119, n28105, n28115, 
        n3_adj_6625, n28111, n22_adj_6626, n28101, n8_adj_6627, n30073, 
        n18610, n10335, n30162, n18456, n26293, n27537, n27545, 
        n27543, n27529, n27539, n3_adj_6628, n27535, n22_adj_6629, 
        n27525, n8_adj_6630, n27513, n27521, n27519, n27505, n27515, 
        n3_adj_6631, n27511, n22_adj_6632, n27501, n8_adj_6633, n27609, 
        n27617, n27615, n27601, n27611, n3_adj_6634, n27607, n22_adj_6635, 
        n27597, n8_adj_6636, n27633, n27641, n27639, n27625, n27635, 
        n3_adj_6637, n27631, n22_adj_6638, n29679, n27621, n8_adj_6639, 
        n27657, n27665, n27663, n27649, n27659, n3_adj_6640, n27655, 
        n22_adj_6641, n27645, n8_adj_6642, n28137, n28145, n28143, 
        n28129, n28139, n3_adj_6643, n28135, n22_adj_6644, n28125, 
        n8_adj_6645, n27921, n27929, n27927, n27913, n27923, n3_adj_6646, 
        n27919, n22_adj_6647, n27909, n8_adj_6648, n27753, n27761, 
        n27759, n27745, n27755, n3_adj_6649, n27751, n22_adj_6650, 
        n27741, n8_adj_6651, n27777, n27785, n27783, n27769, n27779, 
        n3_adj_6652, n27775, n22_adj_6653, n27765, n8_adj_6654, n27897, 
        n27905, n27903, n27889, n27899, n3_adj_6655, n27895, n22_adj_6656, 
        n27885, n8_adj_6657, n27945, n27953, n27951, n27937, n27947, 
        n3_adj_6658, n27943, n22_adj_6659, n27933, n8_adj_6660, n27873, 
        n27881, n27879, n27865, n27875, n3_adj_6661, n27871, n22_adj_6662, 
        n27861, n8_adj_6663, n27993, n28001, n27999, n27985, n27995, 
        n3_adj_6664, n27991, n22_adj_6665, n27981, n8_adj_6666, n29682, 
        n30072, MA_Temp_N_6202, n27705, n27713, n27711, n27697, 
        n27707, n3_adj_6667, n27703, n22_adj_6668, n27693, n8_adj_6669, 
        n28177, n28171, n28173, n22_adj_6670, n28167, n28161, n28163, 
        n22_adj_6671, n28157, n28151, n28153, n22_adj_6672, n30167, 
        n30166, n28187, n28181, n28183, n22_adj_6673, n28197, n28191, 
        n28193, n22_adj_6674, n28207, n28201, n28203, n22_adj_6675, 
        n28217, n28211, n28213, n22_adj_6676, n28227, n28221, n28223, 
        n22_adj_6677, clk_1MHz_enable_57;
    wire [11:0]Cnt_NSL;   // c:/s_links/sources/slot_cards/stepper.v(61[12:19])
    
    wire n30065, n26391, clk_enable_1114, n4, n22086, n22085, n26159, 
        n21974;
    wire [31:0]n153;
    
    wire n22084, n22083, n22082, n22081, n27487, n27497, n27491, 
        n27485, n10_adj_6688, n27469, n27461, n15, n22_adj_6689, 
        n27489, n27481, n8_adj_6690, n27475, n18_adj_6691, n27465, 
        n11_adj_6693, n27477, n5_adj_6696, n30163, n29681, n21973, 
        n21972, n21971, n30192, OW_ID_N_6177, n27447, n27457, n27451, 
        n27445, n27431, n27425, n22_adj_6699, n27449, n27441, n8_adj_6700, 
        n27435, n19_adj_6701, n12588, n27423, n11_adj_6702, n27437, 
        n7_adj_6703, n27825, n27833, n27831, n27817, n27827, n3_adj_6704, 
        n27823, n22_adj_6705, n27813, n8_adj_6706, n27969;
    
    LUT4 i1_4_lut (.A(n27971), .B(\spi_data_out_r_39__N_5540[4] ), .C(n3_c), 
         .D(spi_data_out_r_39__N_5580), .Z(n27977)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut.init = 16'hfefa;
    LUT4 i1_4_lut_adj_310 (.A(\spi_data_out_r_39__N_4511[4] ), .B(n27967), 
         .C(n22_c), .D(spi_data_out_r_39__N_4551), .Z(n27975)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_310.init = 16'hfefc;
    FD1P3AX SLO_buf__i1 (.D(SLO[0]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i1.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_311 (.A(\spi_data_out_r_39__N_1404[4] ), .B(\spi_data_out_r_39__N_1639[4] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27961)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_311.init = 16'heca0;
    LUT4 i1_4_lut_adj_312 (.A(\spi_data_out_r_39__N_1874[4] ), .B(n27957), 
         .C(n8), .D(spi_data_out_r_39__N_1914), .Z(n27971)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_312.init = 16'hfefc;
    LUT4 Select_2910_i3_2_lut (.A(\spi_data_out_r_39__N_1169[4] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_c)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2910_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_313 (.A(\spi_data_out_r_39__N_2109[4] ), .B(\spi_data_out_r_39__N_934[4] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27957)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_313.init = 16'heca0;
    LUT4 Select_2910_i8_2_lut (.A(\spi_data_out_r_39__N_2344[4] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2910_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_314 (.A(\spi_data_out_r_39__N_5197[4] ), .B(\spi_data_out_r_39__N_4854[4] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27967)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_314.init = 16'heca0;
    LUT4 Select_2910_i22_2_lut (.A(spi_data_out_r_39__N_5883[4]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_c)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2910_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_315 (.A(n27681), .B(n27689), .C(n27687), .D(n27673), 
         .Z(\spi_data_out_r[5] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_315.init = 16'hfffe;
    LUT4 i1_4_lut_adj_316 (.A(\spi_data_out_r_39__N_3825[5] ), .B(\spi_data_out_r_39__N_4168[5] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27681)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_316.init = 16'heca0;
    LUT4 i1_4_lut_adj_317 (.A(n27683), .B(\spi_data_out_r_39__N_5540[5] ), 
         .C(n3_adj_6595), .D(spi_data_out_r_39__N_5580), .Z(n27689)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_317.init = 16'hfefa;
    FD1P3IX reset_r_491 (.D(n30028), .SP(clk_enable_46), .CD(n30185), 
            .CK(clk), .Q(reset_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam reset_r_491.GSR = "DISABLED";
    FD1P3AX NSL_484 (.D(NSL_N_6215), .SP(clk_1MHz_enable_9), .CK(clk_1MHz), 
            .Q(NSL)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam NSL_484.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_318 (.A(\spi_data_out_r_39__N_4511[5] ), .B(n27679), 
         .C(n22_adj_6596), .D(spi_data_out_r_39__N_4551), .Z(n27687)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_318.init = 16'hfefc;
    LUT4 i1_4_lut_adj_319 (.A(\spi_data_out_r_39__N_1404[5] ), .B(\spi_data_out_r_39__N_1639[5] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27673)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_319.init = 16'heca0;
    LUT4 i1_4_lut_adj_320 (.A(\spi_data_out_r_39__N_1874[5] ), .B(n27669), 
         .C(n8_adj_6597), .D(spi_data_out_r_39__N_1914), .Z(n27683)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_320.init = 16'hfefc;
    LUT4 Select_2909_i3_2_lut (.A(\spi_data_out_r_39__N_1169[5] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6595)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2909_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_321 (.A(\spi_data_out_r_39__N_2109[5] ), .B(\spi_data_out_r_39__N_934[5] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27669)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_321.init = 16'heca0;
    LUT4 Select_2909_i8_2_lut (.A(\spi_data_out_r_39__N_2344[5] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6597)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2909_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_322 (.A(\spi_data_out_r_39__N_5197[5] ), .B(\spi_data_out_r_39__N_4854[5] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27679)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_322.init = 16'heca0;
    LUT4 Select_2909_i22_2_lut (.A(spi_data_out_r_39__N_5883[5]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6596)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2909_i22_2_lut.init = 16'h8888;
    FD1P3IX mode__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_180), .CD(n30185), 
            .CK(clk), .Q(mode[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i0.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_323 (.A(n28065), .B(n28073), .C(n28071), .D(n28057), 
         .Z(\spi_data_out_r[6] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_323.init = 16'hfffe;
    LUT4 i1_4_lut_adj_324 (.A(\spi_data_out_r_39__N_3825[6] ), .B(\spi_data_out_r_39__N_4168[6] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n28065)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_324.init = 16'heca0;
    LUT4 i1_4_lut_adj_325 (.A(n28067), .B(\spi_data_out_r_39__N_5540[6] ), 
         .C(n3_adj_6598), .D(spi_data_out_r_39__N_5580), .Z(n28073)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_325.init = 16'hfefa;
    LUT4 i1_4_lut_adj_326 (.A(\spi_data_out_r_39__N_4511[6] ), .B(n28063), 
         .C(n22_adj_6599), .D(spi_data_out_r_39__N_4551), .Z(n28071)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_326.init = 16'hfefc;
    LUT4 i1_4_lut_adj_327 (.A(\spi_data_out_r_39__N_1404[6] ), .B(\spi_data_out_r_39__N_1639[6] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n28057)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_327.init = 16'heca0;
    LUT4 i1_4_lut_adj_328 (.A(\spi_data_out_r_39__N_1874[6] ), .B(n28053), 
         .C(n8_adj_6600), .D(spi_data_out_r_39__N_1914), .Z(n28067)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_328.init = 16'hfefc;
    LUT4 Select_2908_i3_2_lut (.A(\spi_data_out_r_39__N_1169[6] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6598)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2908_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_329 (.A(\spi_data_out_r_39__N_2109[6] ), .B(\spi_data_out_r_39__N_934[6] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n28053)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_329.init = 16'heca0;
    LUT4 Select_2908_i8_2_lut (.A(\spi_data_out_r_39__N_2344[6] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6600)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2908_i8_2_lut.init = 16'h8888;
    FD1S3AX prev_MA_Temp_487 (.D(MA_Temp), .CK(clk), .Q(prev_MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam prev_MA_Temp_487.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_330 (.A(\spi_data_out_r_39__N_5197[6] ), .B(\spi_data_out_r_39__N_4854[6] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n28063)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_330.init = 16'heca0;
    LUT4 Select_2908_i22_2_lut (.A(spi_data_out_r_39__N_5883[6]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6599)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2908_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_331 (.A(n27729), .B(n27737), .C(n27735), .D(n27721), 
         .Z(\spi_data_out_r[7] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_331.init = 16'hfffe;
    LUT4 i1_4_lut_adj_332 (.A(\spi_data_out_r_39__N_3825[7] ), .B(\spi_data_out_r_39__N_4168[7] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27729)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_332.init = 16'heca0;
    LUT4 i1_4_lut_adj_333 (.A(n27731), .B(\spi_data_out_r_39__N_5540[7] ), 
         .C(n3_adj_6601), .D(spi_data_out_r_39__N_5580), .Z(n27737)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_333.init = 16'hfefa;
    LUT4 i1_4_lut_adj_334 (.A(\spi_data_out_r_39__N_4511[7] ), .B(n27727), 
         .C(n22_adj_6602), .D(spi_data_out_r_39__N_4551), .Z(n27735)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_334.init = 16'hfefc;
    LUT4 i1_4_lut_adj_335 (.A(\spi_data_out_r_39__N_1404[7] ), .B(\spi_data_out_r_39__N_1639[7] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27721)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_335.init = 16'heca0;
    FD1S3AX prev_MA_489 (.D(n30143), .CK(clk), .Q(prev_MA)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam prev_MA_489.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i0 (.D(spi_data_out_r_39__N_6134[0]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i0.GSR = "DISABLED";
    FD1P3IX Cnt__i0 (.D(n199[0]), .SP(clk_1MHz_enable_49), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i0.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_336 (.A(\spi_data_out_r_39__N_1874[7] ), .B(n27717), 
         .C(n8_adj_6603), .D(spi_data_out_r_39__N_1914), .Z(n27731)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_336.init = 16'hfefc;
    LUT4 Select_2907_i3_2_lut (.A(\spi_data_out_r_39__N_1169[7] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6601)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2907_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_337 (.A(\spi_data_out_r_39__N_2109[7] ), .B(\spi_data_out_r_39__N_934[7] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27717)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_337.init = 16'heca0;
    LUT4 Select_2907_i8_2_lut (.A(\spi_data_out_r_39__N_2344[7] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6603)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2907_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_338 (.A(\spi_data_out_r_39__N_5197[7] ), .B(\spi_data_out_r_39__N_4854[7] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27727)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_338.init = 16'heca0;
    FD1P3AX Cnt_NSL_1784__i0 (.D(n53[0]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784__i0.GSR = "DISABLED";
    LUT4 Select_2907_i22_2_lut (.A(spi_data_out_r_39__N_5883[7]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6602)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2907_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_339 (.A(n27585), .B(n27593), .C(n27591), .D(n27577), 
         .Z(\spi_data_out_r[10] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_339.init = 16'hfffe;
    LUT4 i1_4_lut_adj_340 (.A(\spi_data_out_r_39__N_3825[10] ), .B(\spi_data_out_r_39__N_4168[10] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27585)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_340.init = 16'heca0;
    FD1P3IX mode__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_180), .CD(n30185), 
            .CK(clk), .Q(mode[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i2.GSR = "DISABLED";
    FD1P3IX mode__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_180), .CD(n30185), 
            .CK(clk), .Q(mode[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam mode__i1.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_341 (.A(n27587), .B(\spi_data_out_r_39__N_5540[10] ), 
         .C(n3_adj_6604), .D(spi_data_out_r_39__N_5580), .Z(n27593)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_341.init = 16'hfefa;
    LUT4 i1_4_lut_adj_342 (.A(\spi_data_out_r_39__N_4511[10] ), .B(n27583), 
         .C(n22_adj_6605), .D(spi_data_out_r_39__N_4551), .Z(n27591)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_342.init = 16'hfefc;
    LUT4 i1_4_lut_adj_343 (.A(\spi_data_out_r_39__N_1404[10] ), .B(\spi_data_out_r_39__N_1639[10] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27577)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_343.init = 16'heca0;
    LUT4 i1_4_lut_adj_344 (.A(\spi_data_out_r_39__N_1874[10] ), .B(n27573), 
         .C(n8_adj_6606), .D(spi_data_out_r_39__N_1914), .Z(n27587)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_344.init = 16'hfefc;
    LUT4 Select_2904_i3_2_lut (.A(\spi_data_out_r_39__N_1169[10] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6604)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2904_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_345 (.A(\spi_data_out_r_39__N_2109[10] ), .B(\spi_data_out_r_39__N_934[10] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27573)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_345.init = 16'heca0;
    LUT4 Select_2904_i8_2_lut (.A(\spi_data_out_r_39__N_2344[10] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6606)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2904_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_346 (.A(\spi_data_out_r_39__N_5197[10] ), .B(\spi_data_out_r_39__N_4854[10] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27583)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_346.init = 16'heca0;
    LUT4 Select_2904_i22_2_lut (.A(spi_data_out_r_39__N_5883[10]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6605)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2904_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_347 (.A(n27849), .B(n27857), .C(n27855), .D(n27841), 
         .Z(\spi_data_out_r[11] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_347.init = 16'hfffe;
    LUT4 i1_4_lut_adj_348 (.A(\spi_data_out_r_39__N_3825[11] ), .B(\spi_data_out_r_39__N_4168[11] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27849)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_348.init = 16'heca0;
    LUT4 i1_4_lut_adj_349 (.A(n27851), .B(\spi_data_out_r_39__N_5540[11] ), 
         .C(n3_adj_6607), .D(spi_data_out_r_39__N_5580), .Z(n27857)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_349.init = 16'hfefa;
    LUT4 i1_4_lut_adj_350 (.A(\spi_data_out_r_39__N_4511[11] ), .B(n27847), 
         .C(n22_adj_6608), .D(spi_data_out_r_39__N_4551), .Z(n27855)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_350.init = 16'hfefc;
    LUT4 i1_4_lut_adj_351 (.A(\spi_data_out_r_39__N_1404[11] ), .B(\spi_data_out_r_39__N_1639[11] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27841)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_351.init = 16'heca0;
    LUT4 i1_4_lut_adj_352 (.A(\spi_data_out_r_39__N_1874[11] ), .B(n27837), 
         .C(n8_adj_6609), .D(spi_data_out_r_39__N_1914), .Z(n27851)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_352.init = 16'hfefc;
    LUT4 Select_2903_i3_2_lut (.A(\spi_data_out_r_39__N_1169[11] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6607)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2903_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_353 (.A(\spi_data_out_r_39__N_2109[11] ), .B(\spi_data_out_r_39__N_934[11] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27837)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_353.init = 16'heca0;
    LUT4 Select_2903_i8_2_lut (.A(\spi_data_out_r_39__N_2344[11] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6609)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2903_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_354 (.A(\spi_data_out_r_39__N_5197[11] ), .B(\spi_data_out_r_39__N_4854[11] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27847)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_354.init = 16'heca0;
    LUT4 Select_2903_i22_2_lut (.A(spi_data_out_r_39__N_5883[11]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6608)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2903_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_355 (.A(n28089), .B(n28097), .C(n28095), .D(n28081), 
         .Z(\spi_data_out_r[12] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_355.init = 16'hfffe;
    LUT4 i1_4_lut_adj_356 (.A(\spi_data_out_r_39__N_3825[12] ), .B(\spi_data_out_r_39__N_4168[12] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n28089)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_356.init = 16'heca0;
    LUT4 i1_4_lut_adj_357 (.A(n28091), .B(\spi_data_out_r_39__N_5540[12] ), 
         .C(n3_adj_6610), .D(spi_data_out_r_39__N_5580), .Z(n28097)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_357.init = 16'hfefa;
    LUT4 i1_4_lut_adj_358 (.A(\spi_data_out_r_39__N_4511[12] ), .B(n28087), 
         .C(n22_adj_6611), .D(spi_data_out_r_39__N_4551), .Z(n28095)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_358.init = 16'hfefc;
    LUT4 i1_4_lut_adj_359 (.A(\spi_data_out_r_39__N_1404[12] ), .B(\spi_data_out_r_39__N_1639[12] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n28081)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_359.init = 16'heca0;
    LUT4 i1_4_lut_adj_360 (.A(\spi_data_out_r_39__N_1874[12] ), .B(n28077), 
         .C(n8_adj_6612), .D(spi_data_out_r_39__N_1914), .Z(n28091)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_360.init = 16'hfefc;
    LUT4 Select_2902_i3_2_lut (.A(\spi_data_out_r_39__N_1169[12] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6610)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2902_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_361 (.A(\spi_data_out_r_39__N_2109[12] ), .B(\spi_data_out_r_39__N_934[12] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n28077)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_361.init = 16'heca0;
    LUT4 Select_2902_i8_2_lut (.A(\spi_data_out_r_39__N_2344[12] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6612)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2902_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_362 (.A(\spi_data_out_r_39__N_5197[12] ), .B(\spi_data_out_r_39__N_4854[12] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n28087)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_362.init = 16'heca0;
    LUT4 Select_2902_i22_2_lut (.A(spi_data_out_r_39__N_5883[12]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6611)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2902_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_363 (.A(n27561), .B(n27569), .C(n27567), .D(n27553), 
         .Z(\spi_data_out_r[13] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_363.init = 16'hfffe;
    LUT4 i1_4_lut_adj_364 (.A(\spi_data_out_r_39__N_3825[13] ), .B(\spi_data_out_r_39__N_4168[13] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27561)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_364.init = 16'heca0;
    FD1P3IX digital_output_r_492 (.D(n28550), .SP(clk_enable_222), .CD(n30185), 
            .CK(clk), .Q(digital_output_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(142[8] 164[4])
    defparam digital_output_r_492.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_365 (.A(n27563), .B(\spi_data_out_r_39__N_5540[13] ), 
         .C(n3_adj_6613), .D(spi_data_out_r_39__N_5580), .Z(n27569)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_365.init = 16'hfefa;
    LUT4 i1_4_lut_adj_366 (.A(clk_enable_180), .B(EM_STOP), .C(n25741), 
         .D(n23916), .Z(clk_enable_46)) /* synthesis lut_function=(A+!((C (D))+!B)) */ ;
    defparam i1_4_lut_adj_366.init = 16'haeee;
    LUT4 i1_4_lut_adj_367 (.A(\spi_data_out_r_39__N_4511[13] ), .B(n27559), 
         .C(n22_adj_6614), .D(spi_data_out_r_39__N_4551), .Z(n27567)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_367.init = 16'hfefc;
    LUT4 i1_4_lut_adj_368 (.A(\spi_data_out_r_39__N_1404[13] ), .B(\spi_data_out_r_39__N_1639[13] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27553)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_368.init = 16'heca0;
    LUT4 i1_4_lut_adj_369 (.A(\spi_data_out_r_39__N_1874[13] ), .B(n27549), 
         .C(n8_adj_6615), .D(spi_data_out_r_39__N_1914), .Z(n27563)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_369.init = 16'hfefc;
    LUT4 Select_2901_i3_2_lut (.A(\spi_data_out_r_39__N_1169[13] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6613)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2901_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_370 (.A(\spi_data_out_r_39__N_2109[13] ), .B(\spi_data_out_r_39__N_934[13] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27549)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_370.init = 16'heca0;
    LUT4 Select_2901_i8_2_lut (.A(\spi_data_out_r_39__N_2344[13] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6615)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2901_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_371 (.A(\spi_data_out_r_39__N_5197[13] ), .B(\spi_data_out_r_39__N_4854[13] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27559)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_371.init = 16'heca0;
    LUT4 Select_2901_i22_2_lut (.A(spi_data_out_r_39__N_5883[13]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6614)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2901_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_372 (.A(n28041), .B(n28049), .C(n28047), .D(n28033), 
         .Z(\spi_data_out_r[14] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_372.init = 16'hfffe;
    LUT4 i1_4_lut_adj_373 (.A(\spi_data_out_r_39__N_3825[14] ), .B(\spi_data_out_r_39__N_4168[14] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n28041)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_373.init = 16'heca0;
    LUT4 i1_4_lut_adj_374 (.A(n28043), .B(\spi_data_out_r_39__N_5540[14] ), 
         .C(n3_adj_6616), .D(spi_data_out_r_39__N_5580), .Z(n28049)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_374.init = 16'hfefa;
    LUT4 i1_4_lut_adj_375 (.A(\spi_data_out_r_39__N_4511[14] ), .B(n28039), 
         .C(n22_adj_6617), .D(spi_data_out_r_39__N_4551), .Z(n28047)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_375.init = 16'hfefc;
    LUT4 i1_4_lut_adj_376 (.A(\spi_data_out_r_39__N_1404[14] ), .B(\spi_data_out_r_39__N_1639[14] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n28033)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_376.init = 16'heca0;
    LUT4 i1_4_lut_adj_377 (.A(\spi_data_out_r_39__N_1874[14] ), .B(n28029), 
         .C(n8_adj_6618), .D(spi_data_out_r_39__N_1914), .Z(n28043)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_377.init = 16'hfefc;
    LUT4 Select_2900_i3_2_lut (.A(\spi_data_out_r_39__N_1169[14] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6616)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2900_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_378 (.A(\spi_data_out_r_39__N_2109[14] ), .B(\spi_data_out_r_39__N_934[14] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n28029)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_378.init = 16'heca0;
    LUT4 Select_2900_i8_2_lut (.A(\spi_data_out_r_39__N_2344[14] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6618)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2900_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_379 (.A(\spi_data_out_r_39__N_5197[14] ), .B(\spi_data_out_r_39__N_4854[14] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n28039)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_379.init = 16'heca0;
    LUT4 Select_2900_i22_2_lut (.A(spi_data_out_r_39__N_5883[14]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6617)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2900_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_380 (.A(n27801), .B(n27809), .C(n27807), .D(n27793), 
         .Z(\spi_data_out_r[15] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_380.init = 16'hfffe;
    LUT4 i1_4_lut_adj_381 (.A(\spi_data_out_r_39__N_3825[15] ), .B(\spi_data_out_r_39__N_4168[15] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27801)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_381.init = 16'heca0;
    LUT4 i1_4_lut_adj_382 (.A(n27803), .B(\spi_data_out_r_39__N_5540[15] ), 
         .C(n3_adj_6619), .D(spi_data_out_r_39__N_5580), .Z(n27809)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_382.init = 16'hfefa;
    LUT4 i1_4_lut_adj_383 (.A(\spi_data_out_r_39__N_4511[15] ), .B(n27799), 
         .C(n22_adj_6620), .D(spi_data_out_r_39__N_4551), .Z(n27807)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_383.init = 16'hfefc;
    LUT4 i1_4_lut_adj_384 (.A(\spi_data_out_r_39__N_1404[15] ), .B(\spi_data_out_r_39__N_1639[15] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27793)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_384.init = 16'heca0;
    LUT4 i1_4_lut_adj_385 (.A(\spi_data_out_r_39__N_1874[15] ), .B(n27789), 
         .C(n8_adj_6621), .D(spi_data_out_r_39__N_1914), .Z(n27803)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_385.init = 16'hfefc;
    LUT4 Select_2899_i3_2_lut (.A(\spi_data_out_r_39__N_1169[15] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6619)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2899_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_386 (.A(\spi_data_out_r_39__N_2109[15] ), .B(\spi_data_out_r_39__N_934[15] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27789)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_386.init = 16'heca0;
    LUT4 Select_2899_i8_2_lut (.A(\spi_data_out_r_39__N_2344[15] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6621)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2899_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_387 (.A(\spi_data_out_r_39__N_5197[15] ), .B(\spi_data_out_r_39__N_4854[15] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27799)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_387.init = 16'heca0;
    LUT4 Select_2899_i22_2_lut (.A(spi_data_out_r_39__N_5883[15]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6620)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2899_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_388 (.A(n28017), .B(n28025), .C(n28023), .D(n28009), 
         .Z(\spi_data_out_r[16] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_388.init = 16'hfffe;
    LUT4 i1_4_lut_adj_389 (.A(\spi_data_out_r_39__N_3825[16] ), .B(\spi_data_out_r_39__N_4168[16] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n28017)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_389.init = 16'heca0;
    LUT4 i1_4_lut_adj_390 (.A(n28019), .B(\spi_data_out_r_39__N_5540[16] ), 
         .C(n3_adj_6622), .D(spi_data_out_r_39__N_5580), .Z(n28025)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_390.init = 16'hfefa;
    LUT4 n18534_bdd_4_lut_24559 (.A(n18534), .B(n30164), .C(MA_Temp), 
         .D(Cnt[5]), .Z(n29680)) /* synthesis lut_function=(!(A+(B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam n18534_bdd_4_lut_24559.init = 16'h1450;
    LUT4 i1_4_lut_adj_391 (.A(\spi_data_out_r_39__N_4511[16] ), .B(n28015), 
         .C(n22_adj_6623), .D(spi_data_out_r_39__N_4551), .Z(n28023)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_391.init = 16'hfefc;
    LUT4 i1_4_lut_adj_392 (.A(\spi_data_out_r_39__N_1404[16] ), .B(\spi_data_out_r_39__N_1639[16] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n28009)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_392.init = 16'heca0;
    LUT4 i1_4_lut_adj_393 (.A(\spi_data_out_r_39__N_1874[16] ), .B(n28005), 
         .C(n8_adj_6624), .D(spi_data_out_r_39__N_1914), .Z(n28019)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_393.init = 16'hfefc;
    LUT4 Select_2898_i3_2_lut (.A(\spi_data_out_r_39__N_1169[16] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6622)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2898_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_394 (.A(\spi_data_out_r_39__N_2109[16] ), .B(\spi_data_out_r_39__N_934[16] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n28005)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_394.init = 16'heca0;
    LUT4 Select_2898_i8_2_lut (.A(\spi_data_out_r_39__N_2344[16] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6624)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2898_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_395 (.A(\spi_data_out_r_39__N_5197[16] ), .B(\spi_data_out_r_39__N_4854[16] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n28015)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_395.init = 16'heca0;
    LUT4 Select_2898_i22_2_lut (.A(spi_data_out_r_39__N_5883[16]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6623)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2898_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_396 (.A(n28113), .B(n28121), .C(n28119), .D(n28105), 
         .Z(\spi_data_out_r[17] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_396.init = 16'hfffe;
    LUT4 i1_4_lut_adj_397 (.A(\spi_data_out_r_39__N_3825[17] ), .B(\spi_data_out_r_39__N_4168[17] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n28113)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_397.init = 16'heca0;
    LUT4 i1_4_lut_adj_398 (.A(n28115), .B(\spi_data_out_r_39__N_5540[17] ), 
         .C(n3_adj_6625), .D(spi_data_out_r_39__N_5580), .Z(n28121)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_398.init = 16'hfefa;
    LUT4 i1_4_lut_adj_399 (.A(\spi_data_out_r_39__N_4511[17] ), .B(n28111), 
         .C(n22_adj_6626), .D(spi_data_out_r_39__N_4551), .Z(n28119)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_399.init = 16'hfefc;
    LUT4 i1_4_lut_adj_400 (.A(\spi_data_out_r_39__N_1404[17] ), .B(\spi_data_out_r_39__N_1639[17] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n28105)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_400.init = 16'heca0;
    FD1S3IX i168_494 (.D(spi_data_out_r_39__N_6220), .CK(clk), .CD(n30185), 
            .Q(spi_data_out_r_39__N_5923)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam i168_494.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_401 (.A(\spi_data_out_r_39__N_1874[17] ), .B(n28101), 
         .C(n8_adj_6627), .D(spi_data_out_r_39__N_1914), .Z(n28115)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_401.init = 16'hfefc;
    LUT4 Select_2897_i3_2_lut (.A(\spi_data_out_r_39__N_1169[17] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6625)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2897_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_402 (.A(\spi_data_out_r_39__N_2109[17] ), .B(\spi_data_out_r_39__N_934[17] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n28101)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_402.init = 16'heca0;
    LUT4 Select_2897_i8_2_lut (.A(\spi_data_out_r_39__N_2344[17] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6627)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2897_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_403 (.A(\spi_data_out_r_39__N_5197[17] ), .B(\spi_data_out_r_39__N_4854[17] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n28111)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_403.init = 16'heca0;
    LUT4 i24004_4_lut (.A(NSL), .B(n30073), .C(n18610), .D(n10335), 
         .Z(NSL_N_6215)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C+(D))))) */ ;
    defparam i24004_4_lut.init = 16'h3b37;
    LUT4 i1_4_lut_adj_404 (.A(n30162), .B(n18456), .C(n26293), .D(Cnt[4]), 
         .Z(n18610)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_404.init = 16'hfefa;
    LUT4 Select_2897_i22_2_lut (.A(spi_data_out_r_39__N_5883[17]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6626)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2897_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_405 (.A(n27537), .B(n27545), .C(n27543), .D(n27529), 
         .Z(\spi_data_out_r[18] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_405.init = 16'hfffe;
    LUT4 i1_4_lut_adj_406 (.A(\spi_data_out_r_39__N_3825[18] ), .B(\spi_data_out_r_39__N_4168[18] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27537)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_406.init = 16'heca0;
    LUT4 i1_4_lut_adj_407 (.A(n27539), .B(\spi_data_out_r_39__N_5540[18] ), 
         .C(n3_adj_6628), .D(spi_data_out_r_39__N_5580), .Z(n27545)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_407.init = 16'hfefa;
    LUT4 i1_4_lut_adj_408 (.A(\spi_data_out_r_39__N_4511[18] ), .B(n27535), 
         .C(n22_adj_6629), .D(spi_data_out_r_39__N_4551), .Z(n27543)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_408.init = 16'hfefc;
    LUT4 i1_4_lut_adj_409 (.A(\spi_data_out_r_39__N_1404[18] ), .B(\spi_data_out_r_39__N_1639[18] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27529)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_409.init = 16'heca0;
    LUT4 i1_4_lut_adj_410 (.A(\spi_data_out_r_39__N_1874[18] ), .B(n27525), 
         .C(n8_adj_6630), .D(spi_data_out_r_39__N_1914), .Z(n27539)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_410.init = 16'hfefc;
    LUT4 Select_2896_i3_2_lut (.A(\spi_data_out_r_39__N_1169[18] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6628)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2896_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_411 (.A(\spi_data_out_r_39__N_2109[18] ), .B(\spi_data_out_r_39__N_934[18] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27525)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_411.init = 16'heca0;
    LUT4 Select_2896_i8_2_lut (.A(\spi_data_out_r_39__N_2344[18] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6630)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2896_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_412 (.A(\spi_data_out_r_39__N_5197[18] ), .B(\spi_data_out_r_39__N_4854[18] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27535)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_412.init = 16'heca0;
    LUT4 Select_2896_i22_2_lut (.A(spi_data_out_r_39__N_5883[18]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6629)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2896_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_413 (.A(n27513), .B(n27521), .C(n27519), .D(n27505), 
         .Z(\spi_data_out_r[19] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_413.init = 16'hfffe;
    LUT4 i1_4_lut_adj_414 (.A(\spi_data_out_r_39__N_3825[19] ), .B(\spi_data_out_r_39__N_4168[19] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27513)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_414.init = 16'heca0;
    LUT4 i1_4_lut_adj_415 (.A(n27515), .B(\spi_data_out_r_39__N_5540[19] ), 
         .C(n3_adj_6631), .D(spi_data_out_r_39__N_5580), .Z(n27521)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_415.init = 16'hfefa;
    LUT4 i1_4_lut_adj_416 (.A(\spi_data_out_r_39__N_4511[19] ), .B(n27511), 
         .C(n22_adj_6632), .D(spi_data_out_r_39__N_4551), .Z(n27519)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_416.init = 16'hfefc;
    LUT4 i1_4_lut_adj_417 (.A(\spi_data_out_r_39__N_1404[19] ), .B(\spi_data_out_r_39__N_1639[19] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27505)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_417.init = 16'heca0;
    LUT4 i1_4_lut_adj_418 (.A(\spi_data_out_r_39__N_1874[19] ), .B(n27501), 
         .C(n8_adj_6633), .D(spi_data_out_r_39__N_1914), .Z(n27515)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_418.init = 16'hfefc;
    LUT4 Select_2895_i3_2_lut (.A(\spi_data_out_r_39__N_1169[19] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6631)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2895_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_419 (.A(\spi_data_out_r_39__N_2109[19] ), .B(\spi_data_out_r_39__N_934[19] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27501)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_419.init = 16'heca0;
    LUT4 Select_2895_i8_2_lut (.A(\spi_data_out_r_39__N_2344[19] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6633)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2895_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_420 (.A(\spi_data_out_r_39__N_5197[19] ), .B(\spi_data_out_r_39__N_4854[19] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27511)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_420.init = 16'heca0;
    LUT4 Select_2895_i22_2_lut (.A(spi_data_out_r_39__N_5883[19]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6632)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2895_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_421 (.A(n27609), .B(n27617), .C(n27615), .D(n27601), 
         .Z(\spi_data_out_r[20] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_421.init = 16'hfffe;
    LUT4 i1_4_lut_adj_422 (.A(\spi_data_out_r_39__N_3825[20] ), .B(\spi_data_out_r_39__N_4168[20] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27609)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_422.init = 16'heca0;
    LUT4 i1_4_lut_adj_423 (.A(n27611), .B(\spi_data_out_r_39__N_5540[20] ), 
         .C(n3_adj_6634), .D(spi_data_out_r_39__N_5580), .Z(n27617)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_423.init = 16'hfefa;
    LUT4 i1_4_lut_adj_424 (.A(\spi_data_out_r_39__N_4511[20] ), .B(n27607), 
         .C(n22_adj_6635), .D(spi_data_out_r_39__N_4551), .Z(n27615)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_424.init = 16'hfefc;
    LUT4 i1_4_lut_adj_425 (.A(\spi_data_out_r_39__N_1404[20] ), .B(\spi_data_out_r_39__N_1639[20] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27601)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_425.init = 16'heca0;
    LUT4 i1_4_lut_adj_426 (.A(\spi_data_out_r_39__N_1874[20] ), .B(n27597), 
         .C(n8_adj_6636), .D(spi_data_out_r_39__N_1914), .Z(n27611)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_426.init = 16'hfefc;
    LUT4 Select_2894_i3_2_lut (.A(\spi_data_out_r_39__N_1169[20] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6634)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2894_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_427 (.A(\spi_data_out_r_39__N_2109[20] ), .B(\spi_data_out_r_39__N_934[20] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27597)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_427.init = 16'heca0;
    LUT4 Select_2894_i8_2_lut (.A(\spi_data_out_r_39__N_2344[20] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6636)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2894_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_428 (.A(\spi_data_out_r_39__N_5197[20] ), .B(\spi_data_out_r_39__N_4854[20] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27607)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_428.init = 16'heca0;
    LUT4 Select_2894_i22_2_lut (.A(spi_data_out_r_39__N_5883[20]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6635)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2894_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_429 (.A(n27633), .B(n27641), .C(n27639), .D(n27625), 
         .Z(\spi_data_out_r[21] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_429.init = 16'hfffe;
    LUT4 i1_4_lut_adj_430 (.A(\spi_data_out_r_39__N_3825[21] ), .B(\spi_data_out_r_39__N_4168[21] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27633)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_430.init = 16'heca0;
    LUT4 i1_4_lut_adj_431 (.A(n27635), .B(\spi_data_out_r_39__N_5540[21] ), 
         .C(n3_adj_6637), .D(spi_data_out_r_39__N_5580), .Z(n27641)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_431.init = 16'hfefa;
    LUT4 i1_4_lut_adj_432 (.A(\spi_data_out_r_39__N_4511[21] ), .B(n27631), 
         .C(n22_adj_6638), .D(spi_data_out_r_39__N_4551), .Z(n27639)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_432.init = 16'hfefc;
    LUT4 n18534_bdd_3_lut_24306 (.A(n18534), .B(n18610), .C(MA_Temp), 
         .Z(n29679)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam n18534_bdd_3_lut_24306.init = 16'h7070;
    LUT4 i1_4_lut_adj_433 (.A(\spi_data_out_r_39__N_1404[21] ), .B(\spi_data_out_r_39__N_1639[21] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27625)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_433.init = 16'heca0;
    LUT4 i1_4_lut_adj_434 (.A(\spi_data_out_r_39__N_1874[21] ), .B(n27621), 
         .C(n8_adj_6639), .D(spi_data_out_r_39__N_1914), .Z(n27635)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_434.init = 16'hfefc;
    LUT4 Select_2893_i3_2_lut (.A(\spi_data_out_r_39__N_1169[21] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6637)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2893_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_435 (.A(\spi_data_out_r_39__N_2109[21] ), .B(\spi_data_out_r_39__N_934[21] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27621)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_435.init = 16'heca0;
    LUT4 Select_2893_i8_2_lut (.A(\spi_data_out_r_39__N_2344[21] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6639)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2893_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_436 (.A(\spi_data_out_r_39__N_5197[21] ), .B(\spi_data_out_r_39__N_4854[21] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27631)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_436.init = 16'heca0;
    LUT4 Select_2893_i22_2_lut (.A(spi_data_out_r_39__N_5883[21]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6638)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2893_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_437 (.A(n27657), .B(n27665), .C(n27663), .D(n27649), 
         .Z(\spi_data_out_r[22] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_437.init = 16'hfffe;
    LUT4 i1_4_lut_adj_438 (.A(\spi_data_out_r_39__N_3825[22] ), .B(\spi_data_out_r_39__N_4168[22] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27657)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_438.init = 16'heca0;
    LUT4 i1_4_lut_adj_439 (.A(n27659), .B(\spi_data_out_r_39__N_5540[22] ), 
         .C(n3_adj_6640), .D(spi_data_out_r_39__N_5580), .Z(n27665)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_439.init = 16'hfefa;
    LUT4 i1_4_lut_adj_440 (.A(\spi_data_out_r_39__N_4511[22] ), .B(n27655), 
         .C(n22_adj_6641), .D(spi_data_out_r_39__N_4551), .Z(n27663)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_440.init = 16'hfefc;
    LUT4 i1_4_lut_adj_441 (.A(\spi_data_out_r_39__N_1404[22] ), .B(\spi_data_out_r_39__N_1639[22] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27649)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_441.init = 16'heca0;
    LUT4 i1_4_lut_adj_442 (.A(\spi_data_out_r_39__N_1874[22] ), .B(n27645), 
         .C(n8_adj_6642), .D(spi_data_out_r_39__N_1914), .Z(n27659)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_442.init = 16'hfefc;
    LUT4 Select_2892_i3_2_lut (.A(\spi_data_out_r_39__N_1169[22] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6640)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2892_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_443 (.A(\spi_data_out_r_39__N_2109[22] ), .B(\spi_data_out_r_39__N_934[22] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27645)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_443.init = 16'heca0;
    LUT4 Select_2892_i8_2_lut (.A(\spi_data_out_r_39__N_2344[22] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6642)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2892_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_444 (.A(\spi_data_out_r_39__N_5197[22] ), .B(\spi_data_out_r_39__N_4854[22] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27655)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_444.init = 16'heca0;
    LUT4 Select_2892_i22_2_lut (.A(spi_data_out_r_39__N_5883[22]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6641)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2892_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_445 (.A(n28137), .B(n28145), .C(n28143), .D(n28129), 
         .Z(\spi_data_out_r[23] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_445.init = 16'hfffe;
    LUT4 i1_4_lut_adj_446 (.A(\spi_data_out_r_39__N_3825[23] ), .B(\spi_data_out_r_39__N_4168[23] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n28137)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_446.init = 16'heca0;
    LUT4 i1_4_lut_adj_447 (.A(n28139), .B(\spi_data_out_r_39__N_5540[23] ), 
         .C(n3_adj_6643), .D(spi_data_out_r_39__N_5580), .Z(n28145)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_447.init = 16'hfefa;
    LUT4 i1_4_lut_adj_448 (.A(\spi_data_out_r_39__N_4511[23] ), .B(n28135), 
         .C(n22_adj_6644), .D(spi_data_out_r_39__N_4551), .Z(n28143)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_448.init = 16'hfefc;
    LUT4 i1_4_lut_adj_449 (.A(\spi_data_out_r_39__N_1404[23] ), .B(\spi_data_out_r_39__N_1639[23] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n28129)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_449.init = 16'heca0;
    LUT4 i1_4_lut_adj_450 (.A(\spi_data_out_r_39__N_1874[23] ), .B(n28125), 
         .C(n8_adj_6645), .D(spi_data_out_r_39__N_1914), .Z(n28139)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_450.init = 16'hfefc;
    LUT4 Select_2891_i3_2_lut (.A(\spi_data_out_r_39__N_1169[23] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6643)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2891_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_451 (.A(\spi_data_out_r_39__N_2109[23] ), .B(\spi_data_out_r_39__N_934[23] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n28125)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_451.init = 16'heca0;
    LUT4 Select_2891_i8_2_lut (.A(\spi_data_out_r_39__N_2344[23] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6645)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2891_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_452 (.A(\spi_data_out_r_39__N_5197[23] ), .B(\spi_data_out_r_39__N_4854[23] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n28135)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_452.init = 16'heca0;
    LUT4 Select_2891_i22_2_lut (.A(spi_data_out_r_39__N_5883[23]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6644)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2891_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_453 (.A(n27921), .B(n27929), .C(n27927), .D(n27913), 
         .Z(\spi_data_out_r[24] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_453.init = 16'hfffe;
    LUT4 i1_4_lut_adj_454 (.A(\spi_data_out_r_39__N_3825[24] ), .B(\spi_data_out_r_39__N_4168[24] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27921)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_454.init = 16'heca0;
    LUT4 i1_4_lut_adj_455 (.A(n27923), .B(\spi_data_out_r_39__N_5540[24] ), 
         .C(n3_adj_6646), .D(spi_data_out_r_39__N_5580), .Z(n27929)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_455.init = 16'hfefa;
    LUT4 i1_4_lut_adj_456 (.A(\spi_data_out_r_39__N_4511[24] ), .B(n27919), 
         .C(n22_adj_6647), .D(spi_data_out_r_39__N_4551), .Z(n27927)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_456.init = 16'hfefc;
    LUT4 i1_4_lut_adj_457 (.A(\spi_data_out_r_39__N_1404[24] ), .B(\spi_data_out_r_39__N_1639[24] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27913)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_457.init = 16'heca0;
    LUT4 i1_4_lut_adj_458 (.A(\spi_data_out_r_39__N_1874[24] ), .B(n27909), 
         .C(n8_adj_6648), .D(spi_data_out_r_39__N_1914), .Z(n27923)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_458.init = 16'hfefc;
    LUT4 Select_2890_i3_2_lut (.A(\spi_data_out_r_39__N_1169[24] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6646)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2890_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_459 (.A(\spi_data_out_r_39__N_2109[24] ), .B(\spi_data_out_r_39__N_934[24] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27909)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_459.init = 16'heca0;
    LUT4 Select_2890_i8_2_lut (.A(\spi_data_out_r_39__N_2344[24] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6648)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2890_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_460 (.A(\spi_data_out_r_39__N_5197[24] ), .B(\spi_data_out_r_39__N_4854[24] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27919)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_460.init = 16'heca0;
    LUT4 Select_2890_i22_2_lut (.A(spi_data_out_r_39__N_5883[24]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6647)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2890_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_461 (.A(n27753), .B(n27761), .C(n27759), .D(n27745), 
         .Z(\spi_data_out_r[25] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_461.init = 16'hfffe;
    LUT4 i1_4_lut_adj_462 (.A(\spi_data_out_r_39__N_3825[25] ), .B(\spi_data_out_r_39__N_4168[25] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27753)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_462.init = 16'heca0;
    LUT4 i1_4_lut_adj_463 (.A(n27755), .B(\spi_data_out_r_39__N_5540[25] ), 
         .C(n3_adj_6649), .D(spi_data_out_r_39__N_5580), .Z(n27761)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_463.init = 16'hfefa;
    LUT4 i1_4_lut_adj_464 (.A(\spi_data_out_r_39__N_4511[25] ), .B(n27751), 
         .C(n22_adj_6650), .D(spi_data_out_r_39__N_4551), .Z(n27759)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_464.init = 16'hfefc;
    LUT4 i1_4_lut_adj_465 (.A(\spi_data_out_r_39__N_1404[25] ), .B(\spi_data_out_r_39__N_1639[25] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27745)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_465.init = 16'heca0;
    LUT4 i1_4_lut_adj_466 (.A(\spi_data_out_r_39__N_1874[25] ), .B(n27741), 
         .C(n8_adj_6651), .D(spi_data_out_r_39__N_1914), .Z(n27755)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_466.init = 16'hfefc;
    LUT4 Select_2889_i3_2_lut (.A(\spi_data_out_r_39__N_1169[25] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6649)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2889_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_467 (.A(\spi_data_out_r_39__N_2109[25] ), .B(\spi_data_out_r_39__N_934[25] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27741)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_467.init = 16'heca0;
    LUT4 Select_2889_i8_2_lut (.A(\spi_data_out_r_39__N_2344[25] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6651)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2889_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_468 (.A(\spi_data_out_r_39__N_5197[25] ), .B(\spi_data_out_r_39__N_4854[25] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27751)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_468.init = 16'heca0;
    LUT4 Select_2889_i22_2_lut (.A(spi_data_out_r_39__N_5883[25]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6650)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2889_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_469 (.A(n27777), .B(n27785), .C(n27783), .D(n27769), 
         .Z(\spi_data_out_r[26] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_469.init = 16'hfffe;
    LUT4 i1_4_lut_adj_470 (.A(\spi_data_out_r_39__N_3825[26] ), .B(\spi_data_out_r_39__N_4168[26] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27777)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_470.init = 16'heca0;
    LUT4 i1_4_lut_adj_471 (.A(n27779), .B(\spi_data_out_r_39__N_5540[26] ), 
         .C(n3_adj_6652), .D(spi_data_out_r_39__N_5580), .Z(n27785)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_471.init = 16'hfefa;
    LUT4 i1_4_lut_adj_472 (.A(\spi_data_out_r_39__N_4511[26] ), .B(n27775), 
         .C(n22_adj_6653), .D(spi_data_out_r_39__N_4551), .Z(n27783)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_472.init = 16'hfefc;
    LUT4 i1_4_lut_adj_473 (.A(\spi_data_out_r_39__N_1404[26] ), .B(\spi_data_out_r_39__N_1639[26] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27769)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_473.init = 16'heca0;
    LUT4 i1_4_lut_adj_474 (.A(\spi_data_out_r_39__N_1874[26] ), .B(n27765), 
         .C(n8_adj_6654), .D(spi_data_out_r_39__N_1914), .Z(n27779)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_474.init = 16'hfefc;
    LUT4 Select_2888_i3_2_lut (.A(\spi_data_out_r_39__N_1169[26] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6652)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2888_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_475 (.A(\spi_data_out_r_39__N_2109[26] ), .B(\spi_data_out_r_39__N_934[26] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27765)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_475.init = 16'heca0;
    LUT4 Select_2888_i8_2_lut (.A(\spi_data_out_r_39__N_2344[26] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6654)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2888_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_476 (.A(\spi_data_out_r_39__N_5197[26] ), .B(\spi_data_out_r_39__N_4854[26] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27775)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_476.init = 16'heca0;
    LUT4 Select_2888_i22_2_lut (.A(spi_data_out_r_39__N_5883[26]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6653)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2888_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_477 (.A(n27897), .B(n27905), .C(n27903), .D(n27889), 
         .Z(\spi_data_out_r[27] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_477.init = 16'hfffe;
    LUT4 i1_4_lut_adj_478 (.A(\spi_data_out_r_39__N_3825[27] ), .B(\spi_data_out_r_39__N_4168[27] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27897)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_478.init = 16'heca0;
    LUT4 i1_4_lut_adj_479 (.A(n27899), .B(\spi_data_out_r_39__N_5540[27] ), 
         .C(n3_adj_6655), .D(spi_data_out_r_39__N_5580), .Z(n27905)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_479.init = 16'hfefa;
    LUT4 i1_4_lut_adj_480 (.A(\spi_data_out_r_39__N_4511[27] ), .B(n27895), 
         .C(n22_adj_6656), .D(spi_data_out_r_39__N_4551), .Z(n27903)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_480.init = 16'hfefc;
    LUT4 i1_4_lut_adj_481 (.A(\spi_data_out_r_39__N_1404[27] ), .B(\spi_data_out_r_39__N_1639[27] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27889)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_481.init = 16'heca0;
    LUT4 i1_4_lut_adj_482 (.A(\spi_data_out_r_39__N_1874[27] ), .B(n27885), 
         .C(n8_adj_6657), .D(spi_data_out_r_39__N_1914), .Z(n27899)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_482.init = 16'hfefc;
    LUT4 Select_2887_i3_2_lut (.A(\spi_data_out_r_39__N_1169[27] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6655)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2887_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_483 (.A(\spi_data_out_r_39__N_2109[27] ), .B(\spi_data_out_r_39__N_934[27] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27885)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_483.init = 16'heca0;
    LUT4 Select_2887_i8_2_lut (.A(\spi_data_out_r_39__N_2344[27] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6657)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2887_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_484 (.A(\spi_data_out_r_39__N_5197[27] ), .B(\spi_data_out_r_39__N_4854[27] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27895)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_484.init = 16'heca0;
    LUT4 Select_2887_i22_2_lut (.A(spi_data_out_r_39__N_5883[27]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6656)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2887_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_485 (.A(n27945), .B(n27953), .C(n27951), .D(n27937), 
         .Z(\spi_data_out_r[28] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_485.init = 16'hfffe;
    LUT4 i1_4_lut_adj_486 (.A(\spi_data_out_r_39__N_3825[28] ), .B(\spi_data_out_r_39__N_4168[28] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27945)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_486.init = 16'heca0;
    LUT4 i1_4_lut_adj_487 (.A(n27947), .B(\spi_data_out_r_39__N_5540[28] ), 
         .C(n3_adj_6658), .D(spi_data_out_r_39__N_5580), .Z(n27953)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_487.init = 16'hfefa;
    LUT4 i1_4_lut_adj_488 (.A(\spi_data_out_r_39__N_4511[28] ), .B(n27943), 
         .C(n22_adj_6659), .D(spi_data_out_r_39__N_4551), .Z(n27951)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_488.init = 16'hfefc;
    LUT4 i1_4_lut_adj_489 (.A(\spi_data_out_r_39__N_1404[28] ), .B(\spi_data_out_r_39__N_1639[28] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27937)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_489.init = 16'heca0;
    LUT4 i1_4_lut_adj_490 (.A(\spi_data_out_r_39__N_1874[28] ), .B(n27933), 
         .C(n8_adj_6660), .D(spi_data_out_r_39__N_1914), .Z(n27947)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_490.init = 16'hfefc;
    LUT4 Select_2886_i3_2_lut (.A(\spi_data_out_r_39__N_1169[28] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6658)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2886_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_491 (.A(\spi_data_out_r_39__N_2109[28] ), .B(\spi_data_out_r_39__N_934[28] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27933)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_491.init = 16'heca0;
    LUT4 Select_2886_i8_2_lut (.A(\spi_data_out_r_39__N_2344[28] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6660)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2886_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_492 (.A(\spi_data_out_r_39__N_5197[28] ), .B(\spi_data_out_r_39__N_4854[28] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27943)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_492.init = 16'heca0;
    LUT4 Select_2886_i22_2_lut (.A(spi_data_out_r_39__N_5883[28]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6659)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2886_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_493 (.A(n27873), .B(n27881), .C(n27879), .D(n27865), 
         .Z(\spi_data_out_r[29] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_493.init = 16'hfffe;
    LUT4 i1_4_lut_adj_494 (.A(\spi_data_out_r_39__N_3825[29] ), .B(\spi_data_out_r_39__N_4168[29] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27873)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_494.init = 16'heca0;
    LUT4 i1_4_lut_adj_495 (.A(n27875), .B(\spi_data_out_r_39__N_5540[29] ), 
         .C(n3_adj_6661), .D(spi_data_out_r_39__N_5580), .Z(n27881)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_495.init = 16'hfefa;
    LUT4 i1_4_lut_adj_496 (.A(\spi_data_out_r_39__N_4511[29] ), .B(n27871), 
         .C(n22_adj_6662), .D(spi_data_out_r_39__N_4551), .Z(n27879)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_496.init = 16'hfefc;
    LUT4 i1_4_lut_adj_497 (.A(\spi_data_out_r_39__N_1404[29] ), .B(\spi_data_out_r_39__N_1639[29] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27865)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_497.init = 16'heca0;
    LUT4 i1_4_lut_adj_498 (.A(\spi_data_out_r_39__N_1874[29] ), .B(n27861), 
         .C(n8_adj_6663), .D(spi_data_out_r_39__N_1914), .Z(n27875)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_498.init = 16'hfefc;
    LUT4 Select_2885_i3_2_lut (.A(\spi_data_out_r_39__N_1169[29] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6661)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2885_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_499 (.A(\spi_data_out_r_39__N_2109[29] ), .B(\spi_data_out_r_39__N_934[29] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27861)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_499.init = 16'heca0;
    LUT4 Select_2885_i8_2_lut (.A(\spi_data_out_r_39__N_2344[29] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6663)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2885_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_500 (.A(\spi_data_out_r_39__N_5197[29] ), .B(\spi_data_out_r_39__N_4854[29] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27871)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_500.init = 16'heca0;
    LUT4 i24093_3_lut_4_lut_4_lut (.A(mode[0]), .B(mode[2]), .C(mode[1]), 
         .D(n6), .Z(OW_ID_N_6182)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+!(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(107[27:54])
    defparam i24093_3_lut_4_lut_4_lut.init = 16'hedef;
    LUT4 Select_2885_i22_2_lut (.A(spi_data_out_r_39__N_5883[29]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6662)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2885_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_501 (.A(n27993), .B(n28001), .C(n27999), .D(n27985), 
         .Z(\spi_data_out_r[30] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_501.init = 16'hfffe;
    FD1P3AX SLO_buf__i46 (.D(SLO[45]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i46.GSR = "DISABLED";
    FD1P3AX SLO_buf__i45 (.D(SLO[44]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i45.GSR = "DISABLED";
    FD1P3AX SLO_buf__i44 (.D(SLO[43]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i44.GSR = "DISABLED";
    FD1P3AX SLO_buf__i43 (.D(SLO[42]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i43.GSR = "DISABLED";
    FD1P3AX SLO_buf__i42 (.D(SLO[41]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i42.GSR = "DISABLED";
    FD1P3AX SLO_buf__i41 (.D(SLO[40]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i41.GSR = "DISABLED";
    FD1P3AX SLO_buf__i40 (.D(SLO[39]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i40.GSR = "DISABLED";
    FD1P3AX SLO_buf__i39 (.D(SLO[38]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i39.GSR = "DISABLED";
    FD1P3AX SLO_buf__i38 (.D(SLO[37]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i38.GSR = "DISABLED";
    FD1P3AX SLO_buf__i37 (.D(SLO[36]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i37.GSR = "DISABLED";
    FD1P3AX SLO_buf__i36 (.D(SLO[35]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i36.GSR = "DISABLED";
    FD1P3AX SLO_buf__i35 (.D(SLO[34]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i35.GSR = "DISABLED";
    FD1P3AX SLO_buf__i34 (.D(SLO[33]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i34.GSR = "DISABLED";
    FD1P3AX SLO_buf__i33 (.D(SLO[32]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i33.GSR = "DISABLED";
    FD1P3AX SLO_buf__i32 (.D(SLO[31]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i32.GSR = "DISABLED";
    FD1P3AX SLO_buf__i31 (.D(SLO[30]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i31.GSR = "DISABLED";
    FD1P3AX SLO_buf__i30 (.D(SLO[29]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i30.GSR = "DISABLED";
    FD1P3AX SLO_buf__i29 (.D(SLO[28]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i29.GSR = "DISABLED";
    FD1P3AX SLO_buf__i28 (.D(SLO[27]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i28.GSR = "DISABLED";
    FD1P3AX SLO_buf__i27 (.D(SLO[26]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i27.GSR = "DISABLED";
    FD1P3AX SLO_buf__i26 (.D(SLO[25]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i26.GSR = "DISABLED";
    FD1P3AX SLO_buf__i25 (.D(SLO[24]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i25.GSR = "DISABLED";
    FD1P3AX SLO_buf__i24 (.D(SLO[23]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i24.GSR = "DISABLED";
    FD1P3AX SLO_buf__i23 (.D(SLO[22]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i23.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_502 (.A(\spi_data_out_r_39__N_3825[30] ), .B(\spi_data_out_r_39__N_4168[30] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27993)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_502.init = 16'heca0;
    FD1P3AX SLO_buf__i22 (.D(SLO[21]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i22.GSR = "DISABLED";
    FD1P3AX SLO_buf__i21 (.D(SLO[20]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i21.GSR = "DISABLED";
    FD1P3AX SLO_buf__i20 (.D(SLO[19]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i20.GSR = "DISABLED";
    FD1P3AX SLO_buf__i19 (.D(SLO[18]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i19.GSR = "DISABLED";
    FD1P3AX SLO_buf__i18 (.D(SLO[17]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i18.GSR = "DISABLED";
    FD1P3AX SLO_buf__i17 (.D(SLO[16]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i17.GSR = "DISABLED";
    FD1P3AX SLO_buf__i16 (.D(SLO[15]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i16.GSR = "DISABLED";
    FD1P3AX SLO_buf__i15 (.D(SLO[14]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i15.GSR = "DISABLED";
    FD1P3AX SLO_buf__i14 (.D(SLO[13]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i14.GSR = "DISABLED";
    FD1P3AX SLO_buf__i13 (.D(SLO[12]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i13.GSR = "DISABLED";
    FD1P3AX SLO_buf__i12 (.D(SLO[11]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i12.GSR = "DISABLED";
    FD1P3AX SLO_buf__i11 (.D(SLO[10]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i11.GSR = "DISABLED";
    FD1P3AX SLO_buf__i10 (.D(SLO[9]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i10.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_503 (.A(n27995), .B(\spi_data_out_r_39__N_5540[30] ), 
         .C(n3_adj_6664), .D(spi_data_out_r_39__N_5580), .Z(n28001)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_503.init = 16'hfefa;
    FD1P3AX SLO_buf__i9 (.D(SLO[8]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i9.GSR = "DISABLED";
    FD1P3AX SLO_buf__i8 (.D(SLO[7]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i8.GSR = "DISABLED";
    FD1P3AX SLO_buf__i7 (.D(SLO[6]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i7.GSR = "DISABLED";
    FD1P3AX SLO_buf__i6 (.D(SLO[5]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i6.GSR = "DISABLED";
    FD1P3AX SLO_buf__i5 (.D(SLO[4]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i5.GSR = "DISABLED";
    FD1P3AX SLO_buf__i4 (.D(SLO[3]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i4.GSR = "DISABLED";
    FD1P3AX SLO_buf__i3 (.D(SLO[2]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i3.GSR = "DISABLED";
    FD1P3AX SLO_buf__i2 (.D(SLO[1]), .SP(SLO_buf_51__N_6073), .CK(clk), 
            .Q(SLO_buf[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(121[8] 126[4])
    defparam SLO_buf__i2.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_504 (.A(\spi_data_out_r_39__N_4511[30] ), .B(n27991), 
         .C(n22_adj_6665), .D(spi_data_out_r_39__N_4551), .Z(n27999)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_504.init = 16'hfefc;
    LUT4 i1_4_lut_adj_505 (.A(\spi_data_out_r_39__N_1404[30] ), .B(\spi_data_out_r_39__N_1639[30] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27985)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_505.init = 16'heca0;
    LUT4 i1_4_lut_adj_506 (.A(\spi_data_out_r_39__N_1874[30] ), .B(n27981), 
         .C(n8_adj_6666), .D(spi_data_out_r_39__N_1914), .Z(n27995)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_506.init = 16'hfefc;
    LUT4 n29682_bdd_3_lut (.A(n29682), .B(n29679), .C(n30072), .Z(MA_Temp_N_6202)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n29682_bdd_3_lut.init = 16'hcaca;
    LUT4 Select_2884_i3_2_lut (.A(\spi_data_out_r_39__N_1169[30] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6664)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2884_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_507 (.A(\spi_data_out_r_39__N_2109[30] ), .B(\spi_data_out_r_39__N_934[30] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27981)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_507.init = 16'heca0;
    LUT4 Select_2884_i8_2_lut (.A(\spi_data_out_r_39__N_2344[30] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6666)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2884_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_508 (.A(\spi_data_out_r_39__N_5197[30] ), .B(\spi_data_out_r_39__N_4854[30] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27991)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_508.init = 16'heca0;
    LUT4 Select_2884_i22_2_lut (.A(spi_data_out_r_39__N_5883[30]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6665)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2884_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_509 (.A(n27705), .B(n27713), .C(n27711), .D(n27697), 
         .Z(\spi_data_out_r[31] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_509.init = 16'hfffe;
    LUT4 i1_4_lut_adj_510 (.A(\spi_data_out_r_39__N_3825[31] ), .B(\spi_data_out_r_39__N_4168[31] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27705)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_510.init = 16'heca0;
    LUT4 i1_4_lut_adj_511 (.A(n27707), .B(\spi_data_out_r_39__N_5540[31] ), 
         .C(n3_adj_6667), .D(spi_data_out_r_39__N_5580), .Z(n27713)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_511.init = 16'hfefa;
    LUT4 i1_4_lut_adj_512 (.A(\spi_data_out_r_39__N_4511[31] ), .B(n27703), 
         .C(n22_adj_6668), .D(spi_data_out_r_39__N_4551), .Z(n27711)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_512.init = 16'hfefc;
    LUT4 i1_4_lut_adj_513 (.A(\spi_data_out_r_39__N_1404[31] ), .B(\spi_data_out_r_39__N_1639[31] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27697)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_513.init = 16'heca0;
    LUT4 i1_4_lut_adj_514 (.A(\spi_data_out_r_39__N_1874[31] ), .B(n27693), 
         .C(n8_adj_6669), .D(spi_data_out_r_39__N_1914), .Z(n27707)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_514.init = 16'hfefc;
    LUT4 Select_2883_i3_2_lut (.A(\spi_data_out_r_39__N_1169[31] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6667)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2883_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_515 (.A(\spi_data_out_r_39__N_2109[31] ), .B(\spi_data_out_r_39__N_934[31] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27693)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_515.init = 16'heca0;
    LUT4 Select_2883_i8_2_lut (.A(\spi_data_out_r_39__N_2344[31] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6669)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2883_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_516 (.A(\spi_data_out_r_39__N_5197[31] ), .B(\spi_data_out_r_39__N_4854[31] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27703)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_516.init = 16'heca0;
    LUT4 Select_2883_i22_2_lut (.A(spi_data_out_r_39__N_5883[31]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6668)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2883_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_517 (.A(n28177), .B(n28171), .C(\spi_data_out_r_39__N_4168[32] ), 
         .D(spi_data_out_r_39__N_4208), .Z(\spi_data_out_r[32] )) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_517.init = 16'hfeee;
    LUT4 i1_4_lut_adj_518 (.A(\spi_data_out_r_39__N_4854[32] ), .B(n28173), 
         .C(n22_adj_6670), .D(spi_data_out_r_39__N_4894), .Z(n28177)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_518.init = 16'hfefc;
    LUT4 i1_4_lut_adj_519 (.A(\spi_data_out_r_39__N_5540[32] ), .B(\spi_data_out_r_39__N_4511[32] ), 
         .C(spi_data_out_r_39__N_5580), .D(spi_data_out_r_39__N_4551), .Z(n28171)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_519.init = 16'heca0;
    LUT4 i1_4_lut_adj_520 (.A(\spi_data_out_r_39__N_5197[32] ), .B(\spi_data_out_r_39__N_3825[32] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_3865), .Z(n28173)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_520.init = 16'heca0;
    LUT4 Select_2882_i22_2_lut (.A(spi_data_out_r_39__N_5883[32]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6670)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2882_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_521 (.A(n28167), .B(n28161), .C(\spi_data_out_r_39__N_4168[33] ), 
         .D(spi_data_out_r_39__N_4208), .Z(\spi_data_out_r[33] )) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_521.init = 16'hfeee;
    LUT4 i1_4_lut_adj_522 (.A(\spi_data_out_r_39__N_4854[33] ), .B(n28163), 
         .C(n22_adj_6671), .D(spi_data_out_r_39__N_4894), .Z(n28167)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_522.init = 16'hfefc;
    LUT4 i1_4_lut_adj_523 (.A(\spi_data_out_r_39__N_5540[33] ), .B(\spi_data_out_r_39__N_4511[33] ), 
         .C(spi_data_out_r_39__N_5580), .D(spi_data_out_r_39__N_4551), .Z(n28161)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_523.init = 16'heca0;
    LUT4 i1_4_lut_adj_524 (.A(\spi_data_out_r_39__N_5197[33] ), .B(\spi_data_out_r_39__N_3825[33] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_3865), .Z(n28163)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_524.init = 16'heca0;
    LUT4 Select_2881_i22_2_lut (.A(spi_data_out_r_39__N_5883[33]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6671)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2881_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_525 (.A(n28157), .B(n28151), .C(\spi_data_out_r_39__N_4168[34] ), 
         .D(spi_data_out_r_39__N_4208), .Z(\spi_data_out_r[34] )) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_525.init = 16'hfeee;
    LUT4 i1_4_lut_adj_526 (.A(\spi_data_out_r_39__N_4854[34] ), .B(n28153), 
         .C(n22_adj_6672), .D(spi_data_out_r_39__N_4894), .Z(n28157)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_526.init = 16'hfefc;
    LUT4 i14094_3_lut_4_lut (.A(n30167), .B(n30166), .C(resetn_c), .D(n18610), 
         .Z(clk_1MHz_enable_9)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i14094_3_lut_4_lut.init = 16'h70f0;
    LUT4 i1_4_lut_adj_527 (.A(\spi_data_out_r_39__N_5540[34] ), .B(\spi_data_out_r_39__N_4511[34] ), 
         .C(spi_data_out_r_39__N_5580), .D(spi_data_out_r_39__N_4551), .Z(n28151)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_527.init = 16'heca0;
    LUT4 i1_4_lut_adj_528 (.A(\spi_data_out_r_39__N_5197[34] ), .B(\spi_data_out_r_39__N_3825[34] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_3865), .Z(n28153)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_528.init = 16'heca0;
    LUT4 Select_2880_i22_2_lut (.A(spi_data_out_r_39__N_5883[34]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6672)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2880_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_529 (.A(n28187), .B(n28181), .C(\spi_data_out_r_39__N_4168[35] ), 
         .D(spi_data_out_r_39__N_4208), .Z(\spi_data_out_r[35] )) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_529.init = 16'hfeee;
    LUT4 i1_4_lut_adj_530 (.A(\spi_data_out_r_39__N_4854[35] ), .B(n28183), 
         .C(n22_adj_6673), .D(spi_data_out_r_39__N_4894), .Z(n28187)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_530.init = 16'hfefc;
    LUT4 i1_4_lut_adj_531 (.A(\spi_data_out_r_39__N_5540[35] ), .B(\spi_data_out_r_39__N_4511[35] ), 
         .C(spi_data_out_r_39__N_5580), .D(spi_data_out_r_39__N_4551), .Z(n28181)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_531.init = 16'heca0;
    LUT4 i1_4_lut_adj_532 (.A(\spi_data_out_r_39__N_5197[35] ), .B(\spi_data_out_r_39__N_3825[35] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_3865), .Z(n28183)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_532.init = 16'heca0;
    LUT4 Select_2879_i22_2_lut (.A(spi_data_out_r_39__N_5883[35]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6673)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2879_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_533 (.A(n28197), .B(n28191), .C(\spi_data_out_r_39__N_4168[36] ), 
         .D(spi_data_out_r_39__N_4208), .Z(\spi_data_out_r[36] )) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_533.init = 16'hfeee;
    LUT4 i1_4_lut_adj_534 (.A(\spi_data_out_r_39__N_4854[36] ), .B(n28193), 
         .C(n22_adj_6674), .D(spi_data_out_r_39__N_4894), .Z(n28197)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_534.init = 16'hfefc;
    LUT4 i1_4_lut_adj_535 (.A(\spi_data_out_r_39__N_5540[36] ), .B(\spi_data_out_r_39__N_4511[36] ), 
         .C(spi_data_out_r_39__N_5580), .D(spi_data_out_r_39__N_4551), .Z(n28191)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_535.init = 16'heca0;
    LUT4 i1_4_lut_adj_536 (.A(\spi_data_out_r_39__N_5197[36] ), .B(\spi_data_out_r_39__N_3825[36] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_3865), .Z(n28193)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_536.init = 16'heca0;
    LUT4 Select_2878_i22_2_lut (.A(spi_data_out_r_39__N_5883[36]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6674)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2878_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_537 (.A(n28207), .B(n28201), .C(\spi_data_out_r_39__N_4168[37] ), 
         .D(spi_data_out_r_39__N_4208), .Z(\spi_data_out_r[37] )) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_537.init = 16'hfeee;
    LUT4 i1_4_lut_adj_538 (.A(\spi_data_out_r_39__N_4854[37] ), .B(n28203), 
         .C(n22_adj_6675), .D(spi_data_out_r_39__N_4894), .Z(n28207)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_538.init = 16'hfefc;
    LUT4 i1_4_lut_adj_539 (.A(\spi_data_out_r_39__N_5540[37] ), .B(\spi_data_out_r_39__N_4511[37] ), 
         .C(spi_data_out_r_39__N_5580), .D(spi_data_out_r_39__N_4551), .Z(n28201)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_539.init = 16'heca0;
    LUT4 i1_4_lut_adj_540 (.A(\spi_data_out_r_39__N_5197[37] ), .B(\spi_data_out_r_39__N_3825[37] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_3865), .Z(n28203)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_540.init = 16'heca0;
    LUT4 Select_2877_i22_2_lut (.A(spi_data_out_r_39__N_5883[37]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6675)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2877_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_541 (.A(n28217), .B(n28211), .C(\spi_data_out_r_39__N_4168[38] ), 
         .D(spi_data_out_r_39__N_4208), .Z(\spi_data_out_r[38] )) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_541.init = 16'hfeee;
    LUT4 i1_4_lut_adj_542 (.A(\spi_data_out_r_39__N_4854[38] ), .B(n28213), 
         .C(n22_adj_6676), .D(spi_data_out_r_39__N_4894), .Z(n28217)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_542.init = 16'hfefc;
    LUT4 i1_4_lut_adj_543 (.A(\spi_data_out_r_39__N_5540[38] ), .B(\spi_data_out_r_39__N_4511[38] ), 
         .C(spi_data_out_r_39__N_5580), .D(spi_data_out_r_39__N_4551), .Z(n28211)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_543.init = 16'heca0;
    LUT4 i1_4_lut_adj_544 (.A(\spi_data_out_r_39__N_5197[38] ), .B(\spi_data_out_r_39__N_3825[38] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_3865), .Z(n28213)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_544.init = 16'heca0;
    LUT4 Select_2876_i22_2_lut (.A(spi_data_out_r_39__N_5883[38]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6676)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2876_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_545 (.A(n28227), .B(n28221), .C(\spi_data_out_r_39__N_4168[39] ), 
         .D(spi_data_out_r_39__N_4208), .Z(\spi_data_out_r[39] )) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_545.init = 16'hfeee;
    LUT4 i1_4_lut_adj_546 (.A(\spi_data_out_r_39__N_4854[39] ), .B(n28223), 
         .C(n22_adj_6677), .D(spi_data_out_r_39__N_4894), .Z(n28227)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_546.init = 16'hfefc;
    LUT4 i1_4_lut_adj_547 (.A(\spi_data_out_r_39__N_5540[39] ), .B(\spi_data_out_r_39__N_4511[39] ), 
         .C(spi_data_out_r_39__N_5580), .D(spi_data_out_r_39__N_4551), .Z(n28221)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_547.init = 16'heca0;
    LUT4 i1_4_lut_adj_548 (.A(\spi_data_out_r_39__N_5197[39] ), .B(\spi_data_out_r_39__N_3825[39] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_3865), .Z(n28223)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_548.init = 16'heca0;
    LUT4 Select_2875_i22_2_lut (.A(spi_data_out_r_39__N_5883[39]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6677)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2875_i22_2_lut.init = 16'h8888;
    FD1S3AX spi_data_out_r_i1 (.D(spi_data_out_r_39__N_6134[1]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(spi_data_out_r_39__N_6134[2]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(spi_data_out_r_39__N_6134[3]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(spi_data_out_r_39__N_6134[4]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(spi_data_out_r_39__N_6134[5]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(spi_data_out_r_39__N_6134[6]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(spi_data_out_r_39__N_6134[7]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(spi_data_out_r_39__N_6134[8]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_5883[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(spi_data_out_r_39__N_6134[9]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_5883[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(spi_data_out_r_39__N_6134[10]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(spi_data_out_r_39__N_6134[11]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(spi_data_out_r_39__N_6134[12]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(spi_data_out_r_39__N_6134[13]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(spi_data_out_r_39__N_6134[14]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(spi_data_out_r_39__N_6134[15]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i16 (.D(SLO_buf[30]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i17 (.D(SLO_buf[31]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i18 (.D(SLO_buf[32]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i19 (.D(SLO_buf[33]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i20 (.D(SLO_buf[34]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i21 (.D(SLO_buf[35]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i22 (.D(SLO_buf[36]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i23 (.D(SLO_buf[37]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i24 (.D(SLO_buf[38]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i25 (.D(SLO_buf[39]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i26 (.D(SLO_buf[40]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i27 (.D(SLO_buf[41]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i28 (.D(SLO_buf[42]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i29 (.D(SLO_buf[43]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i30 (.D(SLO_buf[44]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i31 (.D(SLO_buf[45]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(spi_data_out_r_39__N_6134[32]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i33 (.D(spi_data_out_r_39__N_6134[33]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i33.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i34 (.D(spi_data_out_r_39__N_6134[34]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i34.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i35 (.D(spi_data_out_r_39__N_6134[35]), .CK(clk), 
            .Q(spi_data_out_r_39__N_5883[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i35.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i36 (.D(SLO_buf[10]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i36.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i37 (.D(SLO_buf[11]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i37.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i38 (.D(SLO_buf[12]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i38.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i39 (.D(SLO_buf[13]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_5883[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(168[8] 178[4])
    defparam spi_data_out_r_i39.GSR = "DISABLED";
    FD1P3IX Cnt__i1 (.D(n199[1]), .SP(clk_1MHz_enable_49), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i1.GSR = "DISABLED";
    FD1P3IX Cnt__i2 (.D(n199[2]), .SP(clk_1MHz_enable_49), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i3 (.D(n199[3]), .SP(clk_1MHz_enable_49), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i3.GSR = "DISABLED";
    FD1P3IX Cnt__i4 (.D(n199[4]), .SP(clk_1MHz_enable_49), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i4.GSR = "DISABLED";
    FD1P3IX Cnt__i5 (.D(n199[5]), .SP(clk_1MHz_enable_49), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i5.GSR = "DISABLED";
    FD1P3IX Cnt__i6 (.D(n199[6]), .SP(clk_1MHz_enable_49), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i6.GSR = "DISABLED";
    FD1P3IX Cnt__i7 (.D(n199[7]), .SP(clk_1MHz_enable_49), .CD(n30185), 
            .CK(clk_1MHz), .Q(Cnt[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam Cnt__i7.GSR = "DISABLED";
    FD1P3IX MA_Temp_483 (.D(MA_Temp_N_6202), .SP(clk_1MHz_enable_57), .CD(n30185), 
            .CK(clk_1MHz), .Q(MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[8] 115[4])
    defparam MA_Temp_483.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1784__i1 (.D(n53[1]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784__i1.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1784__i2 (.D(n53[2]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784__i2.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1784__i3 (.D(n53[3]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784__i3.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1784__i4 (.D(n53[4]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784__i4.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1784__i5 (.D(n53[5]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784__i5.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1784__i6 (.D(n53[6]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(n93[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784__i6.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1784__i7 (.D(n53[7]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784__i7.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1784__i8 (.D(n53[8]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784__i8.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1784__i9 (.D(n53[9]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784__i9.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1784__i10 (.D(n53[10]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784__i10.GSR = "DISABLED";
    FD1P3AX Cnt_NSL_1784__i11 (.D(n53[11]), .SP(resetn_c), .CK(clk_1MHz), 
            .Q(Cnt_NSL[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784__i11.GSR = "DISABLED";
    LUT4 Select_2906_i16_2_lut (.A(\spi_data_out_r_39__N_3825[8] ), .B(spi_data_out_r_39__N_3865), 
         .Z(n16)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2906_i16_2_lut.init = 16'h8888;
    LUT4 Select_2906_i18_2_lut (.A(\spi_data_out_r_39__N_4511[8] ), .B(spi_data_out_r_39__N_4551), 
         .Z(n18)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2906_i18_2_lut.init = 16'h8888;
    LUT4 Select_2906_i5_2_lut (.A(\spi_data_out_r_39__N_1639[8] ), .B(spi_data_out_r_39__N_1679), 
         .Z(n5)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2906_i5_2_lut.init = 16'h8888;
    LUT4 Select_2906_i3_2_lut (.A(\spi_data_out_r_39__N_1169[8] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2906_i3_2_lut.init = 16'h8888;
    LUT4 Select_2905_i16_2_lut (.A(\spi_data_out_r_39__N_3825[9] ), .B(spi_data_out_r_39__N_3865), 
         .Z(n16_adj_1)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2905_i16_2_lut.init = 16'h8888;
    LUT4 Select_2905_i21_2_lut (.A(\spi_data_out_r_39__N_5540[9] ), .B(spi_data_out_r_39__N_5580), 
         .Z(n21)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2905_i21_2_lut.init = 16'h8888;
    LUT4 Select_2905_i5_2_lut (.A(\spi_data_out_r_39__N_1639[9] ), .B(spi_data_out_r_39__N_1679), 
         .Z(n5_adj_2)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2905_i5_2_lut.init = 16'h8888;
    LUT4 Select_2905_i2_2_lut (.A(\spi_data_out_r_39__N_934[9] ), .B(spi_data_out_r_39__N_974), 
         .Z(n2)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2905_i2_2_lut.init = 16'h8888;
    LUT4 i24144_4_lut (.A(n30065), .B(n26391), .C(n30165), .D(mode[2]), 
         .Z(clk_enable_1114)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C)))) */ ;
    defparam i24144_4_lut.init = 16'h0545;
    LUT4 i1_4_lut_adj_549 (.A(mode[1]), .B(mode[0]), .C(Cnt[4]), .D(n4), 
         .Z(n26391)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut_adj_549.init = 16'h8880;
    LUT4 Select_2912_i21_2_lut (.A(\spi_data_out_r_39__N_5540[2] ), .B(spi_data_out_r_39__N_5580), 
         .Z(n21_adj_3)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2912_i21_2_lut.init = 16'h8888;
    LUT4 Select_2912_i19_2_lut (.A(\spi_data_out_r_39__N_4854[2] ), .B(spi_data_out_r_39__N_4894), 
         .Z(n19)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2912_i19_2_lut.init = 16'h8888;
    CCU2D Cnt_NSL_1784_add_4_13 (.A0(Cnt_NSL[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n22086), .S0(n53[11]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784_add_4_13.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1784_add_4_13.INIT1 = 16'h0000;
    defparam Cnt_NSL_1784_add_4_13.INJECT1_0 = "NO";
    defparam Cnt_NSL_1784_add_4_13.INJECT1_1 = "NO";
    LUT4 Select_2912_i7_2_lut (.A(\spi_data_out_r_39__N_2109[2] ), .B(spi_data_out_r_39__N_2149), 
         .Z(n7)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2912_i7_2_lut.init = 16'h8888;
    CCU2D Cnt_NSL_1784_add_4_11 (.A0(Cnt_NSL[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Cnt_NSL[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22085), .COUT(n22086), .S0(n53[9]), .S1(n53[10]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784_add_4_11.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1784_add_4_11.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1784_add_4_11.INJECT1_0 = "NO";
    defparam Cnt_NSL_1784_add_4_11.INJECT1_1 = "NO";
    LUT4 Select_2912_i22_2_lut (.A(spi_data_out_r_39__N_5883[2]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2912_i22_2_lut.init = 16'h8888;
    LUT4 Select_2912_i14_2_lut (.A(\spi_data_out_r_39__N_2934[2] ), .B(clear_intrpt), 
         .Z(n14)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2912_i14_2_lut.init = 16'h8888;
    LUT4 Select_2912_i9_2_lut (.A(\spi_data_out_r_39__N_2579[2] ), .B(clear_intrpt_adj_4), 
         .Z(n9)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2912_i9_2_lut.init = 16'h8888;
    LUT4 mux_158_i1_3_lut (.A(SLO_buf[14]), .B(SLO_buf[4]), .C(n47), .Z(spi_data_out_r_39__N_6134[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_550 (.A(n26159), .B(Cnt[5]), .C(n18456), .D(Cnt[4]), 
         .Z(n18534)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i1_4_lut_adj_550.init = 16'heaaa;
    CCU2D add_564_9 (.A0(Cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21974), 
          .S0(n153[7]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_9.INIT0 = 16'h5aaa;
    defparam add_564_9.INIT1 = 16'h0000;
    defparam add_564_9.INJECT1_0 = "NO";
    defparam add_564_9.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1784_add_4_9 (.A0(Cnt_NSL[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(Cnt_NSL[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n22084), .COUT(n22085), .S0(n53[7]), .S1(n53[8]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784_add_4_9.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1784_add_4_9.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1784_add_4_9.INJECT1_0 = "NO";
    defparam Cnt_NSL_1784_add_4_9.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1784_add_4_7 (.A0(n93[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n22083), .COUT(n22084), .S0(n53[5]), .S1(n53[6]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784_add_4_7.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1784_add_4_7.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1784_add_4_7.INJECT1_0 = "NO";
    defparam Cnt_NSL_1784_add_4_7.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1784_add_4_5 (.A0(n93[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n22082), .COUT(n22083), .S0(n53[3]), .S1(n53[4]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784_add_4_5.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1784_add_4_5.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1784_add_4_5.INJECT1_0 = "NO";
    defparam Cnt_NSL_1784_add_4_5.INJECT1_1 = "NO";
    CCU2D Cnt_NSL_1784_add_4_3 (.A0(n93[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n93[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n22081), .COUT(n22082), .S0(n53[1]), .S1(n53[2]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784_add_4_3.INIT0 = 16'hfaaa;
    defparam Cnt_NSL_1784_add_4_3.INIT1 = 16'hfaaa;
    defparam Cnt_NSL_1784_add_4_3.INJECT1_0 = "NO";
    defparam Cnt_NSL_1784_add_4_3.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_762 (.A(Cnt[7]), .B(Cnt[6]), .Z(n30162)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(109[8:17])
    defparam i1_2_lut_rep_762.init = 16'heeee;
    LUT4 i1_4_lut_adj_551 (.A(n27487), .B(n27497), .C(n27491), .D(n27485), 
         .Z(\spi_data_out_r[0] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_551.init = 16'hfffe;
    LUT4 i1_4_lut_adj_552 (.A(n10_adj_6688), .B(n27469), .C(n27461), .D(n15), 
         .Z(n27487)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_552.init = 16'hfffe;
    LUT4 i1_4_lut_adj_553 (.A(n22_adj_6689), .B(n27489), .C(n27481), .D(n8_adj_6690), 
         .Z(n27497)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_553.init = 16'hfffe;
    LUT4 i1_4_lut_adj_554 (.A(\spi_data_out_r_39__N_4854[0] ), .B(n27475), 
         .C(n18_adj_6691), .D(spi_data_out_r_39__N_4894), .Z(n27491)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_554.init = 16'hfefc;
    LUT4 i1_4_lut_adj_555 (.A(\spi_data_out_r_39__N_4168[0] ), .B(\spi_data_out_r_39__N_5197[0] ), 
         .C(spi_data_out_r_39__N_4208), .D(spi_data_out_r_39__N_5237), .Z(n27485)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_555.init = 16'heca0;
    LUT4 Select_2914_i10_2_lut (.A(\spi_data_out_r_39__N_2650[0] ), .B(clear_intrpt_adj_5), 
         .Z(n10_adj_6688)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2914_i10_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_556 (.A(\spi_data_out_r_39__N_2863[0] ), .B(n27465), 
         .C(n11_adj_6693), .D(clear_intrpt_adj_6), .Z(n27469)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_556.init = 16'hfefc;
    LUT4 i1_4_lut_adj_557 (.A(\spi_data_out_r_39__N_2934[0] ), .B(\spi_data_out_r_39__N_770[0] ), 
         .C(clear_intrpt), .D(spi_data_out_r_39__N_810), .Z(n27461)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_557.init = 16'heca0;
    LUT4 Select_2914_i15_2_lut (.A(\spi_data_out_r_39__N_3005[0] ), .B(clear_intrpt_adj_7), 
         .Z(n15)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2914_i15_2_lut.init = 16'h8888;
    LUT4 Select_2914_i22_2_lut (.A(spi_data_out_r_39__N_5883[0]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6689)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2914_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_558 (.A(\spi_data_out_r_39__N_2109[0] ), .B(n27477), 
         .C(n5_adj_6696), .D(spi_data_out_r_39__N_2149), .Z(n27489)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_558.init = 16'hfefc;
    LUT4 i1_4_lut_adj_559 (.A(\spi_data_out_r_39__N_3825[0] ), .B(\spi_data_out_r_39__N_5540[0] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_5580), .Z(n27481)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_559.init = 16'heca0;
    LUT4 Select_2914_i8_2_lut (.A(\spi_data_out_r_39__N_2344[0] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6690)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2914_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_560 (.A(\spi_data_out_r_39__N_934[0] ), .B(\spi_data_out_r_39__N_1404[0] ), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_1444), .Z(n27477)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_560.init = 16'heca0;
    LUT4 Select_2914_i5_2_lut (.A(\spi_data_out_r_39__N_1639[0] ), .B(spi_data_out_r_39__N_1679), 
         .Z(n5_adj_6696)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2914_i5_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_561 (.A(\spi_data_out_r_39__N_1169[0] ), .B(\spi_data_out_r_39__N_1874[0] ), 
         .C(spi_data_out_r_39__N_1209), .D(spi_data_out_r_39__N_1914), .Z(n27475)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_561.init = 16'heca0;
    LUT4 Select_2914_i18_2_lut (.A(\spi_data_out_r_39__N_4511[0] ), .B(spi_data_out_r_39__N_4551), 
         .Z(n18_adj_6691)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2914_i18_2_lut.init = 16'h8888;
    CCU2D Cnt_NSL_1784_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n30166), .B1(n30167), .C1(n93[0]), .D1(GND_net), 
          .COUT(n22081), .S1(n53[0]));   // c:/s_links/sources/slot_cards/stepper.v(100[15:26])
    defparam Cnt_NSL_1784_add_4_1.INIT0 = 16'hF000;
    defparam Cnt_NSL_1784_add_4_1.INIT1 = 16'h8787;
    defparam Cnt_NSL_1784_add_4_1.INJECT1_0 = "NO";
    defparam Cnt_NSL_1784_add_4_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_562 (.A(\spi_data_out_r_39__N_2792[0] ), .B(\spi_data_out_r_39__N_2579[0] ), 
         .C(clear_intrpt_adj_8), .D(clear_intrpt_adj_4), .Z(n27465)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_562.init = 16'heca0;
    LUT4 Select_2914_i11_2_lut (.A(\spi_data_out_r_39__N_2721[0] ), .B(clear_intrpt_adj_9), 
         .Z(n11_adj_6693)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2914_i11_2_lut.init = 16'h8888;
    LUT4 i1_3_lut_rep_672_4_lut (.A(Cnt[7]), .B(Cnt[6]), .C(Cnt[0]), .D(n30163), 
         .Z(n30072)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(109[8:17])
    defparam i1_3_lut_rep_672_4_lut.init = 16'hfffe;
    PFUMX i24307 (.BLUT(n29681), .ALUT(n29680), .C0(n18610), .Z(n29682));
    CCU2D add_564_7 (.A0(Cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21973), 
          .COUT(n21974), .S0(n153[5]), .S1(n153[6]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_7.INIT0 = 16'h5aaa;
    defparam add_564_7.INIT1 = 16'h5aaa;
    defparam add_564_7.INJECT1_0 = "NO";
    defparam add_564_7.INJECT1_1 = "NO";
    CCU2D add_564_5 (.A0(Cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21972), 
          .COUT(n21973), .S0(n153[3]), .S1(n153[4]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_5.INIT0 = 16'h5aaa;
    defparam add_564_5.INIT1 = 16'h5aaa;
    defparam add_564_5.INJECT1_0 = "NO";
    defparam add_564_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_763 (.A(Cnt[2]), .B(Cnt[3]), .Z(n30163)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(109[8:17])
    defparam i1_2_lut_rep_763.init = 16'heeee;
    LUT4 i1_3_lut_4_lut (.A(Cnt[2]), .B(Cnt[3]), .C(Cnt[1]), .D(Cnt[0]), 
         .Z(n18456)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(109[8:17])
    defparam i1_3_lut_4_lut.init = 16'hfeee;
    LUT4 i13285_2_lut_rep_764 (.A(Cnt[4]), .B(Cnt[1]), .Z(n30164)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13285_2_lut_rep_764.init = 16'h8888;
    LUT4 n18534_bdd_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(Cnt[5]), .D(MA_Temp), 
         .Z(n29681)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;
    defparam n18534_bdd_3_lut_4_lut.init = 16'hf708;
    LUT4 i1_2_lut_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(n30072), .D(Cnt[5]), 
         .Z(n10335)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff7;
    LUT4 i1_3_lut_rep_765 (.A(mode[1]), .B(mode[2]), .C(mode[0]), .Z(n30165)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_3_lut_rep_765.init = 16'hfbfb;
    CCU2D add_564_3 (.A0(Cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n21971), 
          .COUT(n21972), .S0(n153[1]), .S1(n153[2]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_3.INIT0 = 16'h5aaa;
    defparam add_564_3.INIT1 = 16'h5aaa;
    defparam add_564_3.INJECT1_0 = "NO";
    defparam add_564_3.INJECT1_1 = "NO";
    CCU2D add_564_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n21971), 
          .S1(n153[0]));   // c:/s_links/sources/slot_cards/stepper.v(108[11:16])
    defparam add_564_1.INIT0 = 16'hF000;
    defparam add_564_1.INIT1 = 16'h5555;
    defparam add_564_1.INJECT1_0 = "NO";
    defparam add_564_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(mode[1]), .B(mode[2]), .C(mode[0]), .D(Cnt[5]), 
         .Z(n26293)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i1_2_lut_4_lut.init = 16'hfffb;
    LUT4 i2_3_lut_4_lut (.A(mode[1]), .B(n30192), .C(\uart_slot_en[3] ), 
         .D(pin_io_out_65), .Z(n24700)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(70[15:39])
    defparam i2_3_lut_4_lut.init = 16'he000;
    LUT4 i1_3_lut_rep_766 (.A(Cnt_NSL[9]), .B(Cnt_NSL[8]), .C(Cnt_NSL[7]), 
         .Z(n30166)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_rep_766.init = 16'hfefe;
    LUT4 i1_2_lut_rep_673_4_lut (.A(Cnt_NSL[9]), .B(Cnt_NSL[8]), .C(Cnt_NSL[7]), 
         .D(n30167), .Z(n30073)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_rep_673_4_lut.init = 16'hfe00;
    LUT4 i1_2_lut_rep_767 (.A(Cnt_NSL[11]), .B(Cnt_NSL[10]), .Z(n30167)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i1_2_lut_rep_767.init = 16'h8888;
    LUT4 i23934_2_lut_rep_624_3_lut_4_lut (.A(Cnt_NSL[11]), .B(Cnt_NSL[10]), 
         .C(resetn_c), .D(n30166), .Z(clk_1MHz_enable_49)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(C)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(98[15:29])
    defparam i23934_2_lut_rep_624_3_lut_4_lut.init = 16'h8f0f;
    LUT4 i13013_2_lut_3_lut (.A(n18534), .B(n18610), .C(n153[0]), .Z(n199[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13013_2_lut_3_lut.init = 16'h7070;
    LUT4 i13640_2_lut_3_lut (.A(n18534), .B(n18610), .C(n153[1]), .Z(n199[1])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13640_2_lut_3_lut.init = 16'h7070;
    LUT4 i13641_2_lut_3_lut (.A(n18534), .B(n18610), .C(n153[2]), .Z(n199[2])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13641_2_lut_3_lut.init = 16'h7070;
    LUT4 i13642_2_lut_3_lut (.A(n18534), .B(n18610), .C(n153[3]), .Z(n199[3])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13642_2_lut_3_lut.init = 16'h7070;
    LUT4 i13643_2_lut_3_lut (.A(n18534), .B(n18610), .C(n153[4]), .Z(n199[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13643_2_lut_3_lut.init = 16'h7070;
    LUT4 i13644_2_lut_3_lut (.A(n18534), .B(n18610), .C(n153[5]), .Z(n199[5])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13644_2_lut_3_lut.init = 16'h7070;
    LUT4 i13645_2_lut_3_lut (.A(n18534), .B(n18610), .C(n153[6]), .Z(n199[6])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13645_2_lut_3_lut.init = 16'h7070;
    LUT4 i13646_2_lut_3_lut (.A(n18534), .B(n18610), .C(n153[7]), .Z(n199[7])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13646_2_lut_3_lut.init = 16'h7070;
    LUT4 i2997_2_lut_4_lut (.A(mode[1]), .B(mode[0]), .C(mode[2]), .D(pin_io_c_68), 
         .Z(\quad_a[6] )) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i2997_2_lut_4_lut.init = 16'h0400;
    LUT4 i2998_2_lut_4_lut (.A(mode[1]), .B(mode[0]), .C(mode[2]), .D(pin_io_out_69), 
         .Z(\quad_b[6] )) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[17:38])
    defparam i2998_2_lut_4_lut.init = 16'h0400;
    LUT4 mux_158_i2_3_lut (.A(SLO_buf[15]), .B(SLO_buf[5]), .C(n47), .Z(spi_data_out_r_39__N_6134[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i2_3_lut.init = 16'hcaca;
    LUT4 mux_158_i3_3_lut (.A(SLO_buf[16]), .B(SLO_buf[6]), .C(n47), .Z(spi_data_out_r_39__N_6134[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i3_3_lut.init = 16'hcaca;
    LUT4 mux_158_i4_3_lut (.A(SLO_buf[17]), .B(SLO_buf[7]), .C(n47), .Z(spi_data_out_r_39__N_6134[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i4_3_lut.init = 16'hcaca;
    LUT4 mux_158_i5_3_lut (.A(SLO_buf[18]), .B(SLO_buf[8]), .C(n47), .Z(spi_data_out_r_39__N_6134[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i5_3_lut.init = 16'hcaca;
    LUT4 mux_158_i6_3_lut (.A(SLO_buf[19]), .B(SLO_buf[9]), .C(n47), .Z(spi_data_out_r_39__N_6134[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i6_3_lut.init = 16'hcaca;
    LUT4 mux_158_i7_3_lut (.A(SLO_buf[20]), .B(SLO_buf[10]), .C(n47), 
         .Z(spi_data_out_r_39__N_6134[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i7_3_lut.init = 16'hcaca;
    LUT4 mux_158_i8_3_lut (.A(SLO_buf[21]), .B(SLO_buf[11]), .C(n47), 
         .Z(spi_data_out_r_39__N_6134[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i8_3_lut.init = 16'hcaca;
    LUT4 mux_158_i9_3_lut (.A(SLO_buf[22]), .B(SLO_buf[12]), .C(n47), 
         .Z(spi_data_out_r_39__N_6134[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i9_3_lut.init = 16'hcaca;
    LUT4 digital_output_r_I_0_547_3_lut (.A(digital_output_r), .B(UC_TXD0_c), 
         .C(OW_ID_N_6177), .Z(OW_ID_N_6176)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(90[16] 91[59])
    defparam digital_output_r_I_0_547_3_lut.init = 16'hcaca;
    LUT4 mux_158_i10_3_lut (.A(SLO_buf[23]), .B(SLO_buf[13]), .C(n47), 
         .Z(spi_data_out_r_39__N_6134[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i10_3_lut.init = 16'hcaca;
    LUT4 mux_158_i11_3_lut (.A(SLO_buf[24]), .B(SLO_buf[14]), .C(n47), 
         .Z(spi_data_out_r_39__N_6134[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i11_3_lut.init = 16'hcaca;
    LUT4 i4_4_lut (.A(mode[0]), .B(mode[2]), .C(mode[1]), .D(n6), .Z(OW_ID_N_6177)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i4_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_rep_792 (.A(mode[0]), .B(mode[2]), .Z(n30192)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(107[27:54])
    defparam i1_2_lut_rep_792.init = 16'heeee;
    LUT4 i1_2_lut_rep_683_3_lut (.A(mode[0]), .B(mode[2]), .C(mode[1]), 
         .Z(n30083)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(107[27:54])
    defparam i1_2_lut_rep_683_3_lut.init = 16'hfefe;
    LUT4 i2995_2_lut_3_lut_4_lut (.A(mode[0]), .B(mode[2]), .C(pin_io_c_63), 
         .D(mode[1]), .Z(\pin_intrpt[19] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(107[27:54])
    defparam i2995_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2996_2_lut_3_lut_4_lut (.A(mode[0]), .B(mode[2]), .C(pin_io_c_64), 
         .D(mode[1]), .Z(\pin_intrpt[20] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(107[27:54])
    defparam i2996_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2994_2_lut_3_lut_4_lut (.A(mode[0]), .B(mode[2]), .C(pin_io_c_62), 
         .D(mode[1]), .Z(\pin_intrpt[18] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(107[27:54])
    defparam i2994_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2944_1_lut_2_lut_3_lut (.A(mode[0]), .B(mode[2]), .C(mode[1]), 
         .Z(n7258)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(107[27:54])
    defparam i2944_1_lut_2_lut_3_lut.init = 16'h0101;
    LUT4 mux_158_i12_3_lut (.A(SLO_buf[25]), .B(SLO_buf[15]), .C(n47), 
         .Z(spi_data_out_r_39__N_6134[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i12_3_lut.init = 16'hcaca;
    LUT4 mux_158_i13_3_lut (.A(SLO_buf[26]), .B(SLO_buf[16]), .C(n47), 
         .Z(spi_data_out_r_39__N_6134[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i13_3_lut.init = 16'hcaca;
    LUT4 mux_158_i14_3_lut (.A(SLO_buf[27]), .B(SLO_buf[17]), .C(n47), 
         .Z(spi_data_out_r_39__N_6134[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i14_3_lut.init = 16'hcaca;
    LUT4 mux_158_i15_3_lut (.A(SLO_buf[28]), .B(SLO_buf[18]), .C(n47), 
         .Z(spi_data_out_r_39__N_6134[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i15_3_lut.init = 16'hcaca;
    LUT4 mux_158_i16_3_lut (.A(SLO_buf[29]), .B(SLO_buf[19]), .C(n47), 
         .Z(spi_data_out_r_39__N_6134[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i16_3_lut.init = 16'hcaca;
    LUT4 mux_158_i33_3_lut (.A(SLO_buf[6]), .B(SLO_buf[0]), .C(n47), .Z(spi_data_out_r_39__N_6134[32])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i33_3_lut.init = 16'hcaca;
    LUT4 mux_158_i34_3_lut (.A(SLO_buf[7]), .B(SLO_buf[1]), .C(n47), .Z(spi_data_out_r_39__N_6134[33])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i34_3_lut.init = 16'hcaca;
    LUT4 mux_158_i35_3_lut (.A(SLO_buf[8]), .B(SLO_buf[2]), .C(n47), .Z(spi_data_out_r_39__N_6134[34])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i35_3_lut.init = 16'hcaca;
    LUT4 mux_158_i36_3_lut (.A(SLO_buf[9]), .B(SLO_buf[3]), .C(n47), .Z(spi_data_out_r_39__N_6134[35])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(173[11] 177[5])
    defparam mux_158_i36_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(\quad_homing[0] ), .B(pin_io_c_64), .Z(n25889)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(74[8:17])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i23998_2_lut_3_lut_4_lut (.A(resetn_c), .B(n30073), .C(n18610), 
         .D(n18534), .Z(clk_1MHz_enable_57)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (C (D)))) */ ;
    defparam i23998_2_lut_3_lut_4_lut.init = 16'h0ddd;
    LUT4 i1_4_lut_adj_563 (.A(n27447), .B(n27457), .C(n27451), .D(n27445), 
         .Z(\spi_data_out_r[1] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_563.init = 16'hfffe;
    LUT4 i1_4_lut_adj_564 (.A(n27431), .B(n27425), .C(\spi_data_out_r_39__N_2934[1] ), 
         .D(clear_intrpt), .Z(n27447)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_564.init = 16'hfeee;
    LUT4 i1_4_lut_adj_565 (.A(n22_adj_6699), .B(n27449), .C(n27441), .D(n8_adj_6700), 
         .Z(n27457)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_565.init = 16'hfffe;
    LUT4 i1_4_lut_adj_566 (.A(\spi_data_out_r_39__N_4511[1] ), .B(n27435), 
         .C(n19_adj_6701), .D(spi_data_out_r_39__N_4551), .Z(n27451)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_566.init = 16'hfefc;
    LUT4 i1_4_lut_adj_567 (.A(\spi_data_out_r_39__N_5197[1] ), .B(\spi_data_out_r_39__N_3825[1] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_3865), .Z(n27445)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_567.init = 16'heca0;
    FD1P3IX SLO__i45 (.D(SLO[43]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i45.GSR = "DISABLED";
    FD1P3IX SLO__i46 (.D(SLO[44]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i46.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_568 (.A(\spi_data_out_r_39__N_2863[1] ), .B(n27423), 
         .C(n11_adj_6702), .D(clear_intrpt_adj_6), .Z(n27431)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_568.init = 16'hfefc;
    LUT4 i1_4_lut_adj_569 (.A(\spi_data_out_r_39__N_3005[1] ), .B(\spi_data_out_r_39__N_2579[1] ), 
         .C(clear_intrpt_adj_7), .D(clear_intrpt_adj_4), .Z(n27425)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_569.init = 16'heca0;
    LUT4 i1_4_lut_adj_570 (.A(\spi_data_out_r_39__N_2792[1] ), .B(\spi_data_out_r_39__N_2650[1] ), 
         .C(clear_intrpt_adj_8), .D(clear_intrpt_adj_5), .Z(n27423)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_570.init = 16'heca0;
    LUT4 Select_2913_i11_2_lut (.A(\spi_data_out_r_39__N_2721[1] ), .B(clear_intrpt_adj_9), 
         .Z(n11_adj_6702)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2913_i11_2_lut.init = 16'h8888;
    FD1P3IX SLO__i35 (.D(SLO[33]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i35.GSR = "DISABLED";
    FD1P3IX SLO__i39 (.D(SLO[37]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i39.GSR = "DISABLED";
    FD1P3IX SLO__i42 (.D(SLO[40]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i42.GSR = "DISABLED";
    FD1P3IX SLO__i36 (.D(SLO[34]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i36.GSR = "DISABLED";
    FD1P3IX SLO__i40 (.D(SLO[38]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i40.GSR = "DISABLED";
    FD1P3IX SLO__i43 (.D(SLO[41]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i43.GSR = "DISABLED";
    FD1P3IX SLO__i33 (.D(SLO[31]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i33.GSR = "DISABLED";
    FD1P3IX SLO__i37 (.D(SLO[35]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i37.GSR = "DISABLED";
    FD1P3IX SLO__i34 (.D(SLO[32]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i34.GSR = "DISABLED";
    FD1P3IX SLO__i38 (.D(SLO[36]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i38.GSR = "DISABLED";
    FD1P3IX SLO__i41 (.D(SLO[39]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i41.GSR = "DISABLED";
    FD1P3IX SLO__i44 (.D(SLO[42]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i44.GSR = "DISABLED";
    LUT4 Select_2913_i22_2_lut (.A(spi_data_out_r_39__N_5883[1]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6699)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2913_i22_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_571 (.A(\spi_data_out_r_39__N_1169[1] ), .B(n27437), 
         .C(n7_adj_6703), .D(spi_data_out_r_39__N_1209), .Z(n27449)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_571.init = 16'hfefc;
    LUT4 i1_4_lut_adj_572 (.A(\spi_data_out_r_39__N_4168[1] ), .B(\spi_data_out_r_39__N_5540[1] ), 
         .C(spi_data_out_r_39__N_4208), .D(spi_data_out_r_39__N_5580), .Z(n27441)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_572.init = 16'heca0;
    LUT4 Select_2913_i8_2_lut (.A(\spi_data_out_r_39__N_2344[1] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6700)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2913_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_573 (.A(\spi_data_out_r_39__N_1639[1] ), .B(\spi_data_out_r_39__N_934[1] ), 
         .C(spi_data_out_r_39__N_1679), .D(spi_data_out_r_39__N_974), .Z(n27437)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_573.init = 16'heca0;
    LUT4 Select_2913_i7_2_lut (.A(\spi_data_out_r_39__N_2109[1] ), .B(spi_data_out_r_39__N_2149), 
         .Z(n7_adj_6703)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2913_i7_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_574 (.A(\spi_data_out_r_39__N_1404[1] ), .B(\spi_data_out_r_39__N_1874[1] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1914), .Z(n27435)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_574.init = 16'heca0;
    LUT4 Select_2913_i19_2_lut (.A(\spi_data_out_r_39__N_4854[1] ), .B(spi_data_out_r_39__N_4894), 
         .Z(n19_adj_6701)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2913_i19_2_lut.init = 16'h8888;
    FD1P3IX SLO__i23 (.D(SLO[21]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i23.GSR = "DISABLED";
    FD1P3IX SLO__i27 (.D(SLO[25]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i27.GSR = "DISABLED";
    FD1P3IX SLO__i30 (.D(SLO[28]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i30.GSR = "DISABLED";
    FD1P3IX SLO__i24 (.D(SLO[22]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i24.GSR = "DISABLED";
    FD1P3IX SLO__i28 (.D(SLO[26]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i28.GSR = "DISABLED";
    FD1P3IX SLO__i31 (.D(SLO[29]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i31.GSR = "DISABLED";
    FD1P3IX SLO__i21 (.D(SLO[19]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i21.GSR = "DISABLED";
    FD1P3IX SLO__i25 (.D(SLO[23]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i25.GSR = "DISABLED";
    FD1P3IX SLO__i22 (.D(SLO[20]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i22.GSR = "DISABLED";
    FD1P3IX SLO__i26 (.D(SLO[24]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i26.GSR = "DISABLED";
    FD1P3IX SLO__i29 (.D(SLO[27]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i29.GSR = "DISABLED";
    FD1P3IX SLO__i32 (.D(SLO[30]), .SP(clk_enable_1114), .CD(n12588), 
            .CK(clk), .Q(SLO[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i32.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut (.A(Cnt[5]), .B(n30072), .C(Cnt[1]), .Z(n4)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(133[16:19])
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_575 (.A(n27825), .B(n27833), .C(n27831), .D(n27817), 
         .Z(\spi_data_out_r[3] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_575.init = 16'hfffe;
    LUT4 i1_4_lut_adj_576 (.A(\spi_data_out_r_39__N_3825[3] ), .B(\spi_data_out_r_39__N_4168[3] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27825)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_576.init = 16'heca0;
    FD1P3IX SLO__i12 (.D(SLO[10]), .SP(clk_enable_1114), .CD(GND_net), 
            .CK(clk), .Q(SLO[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i12.GSR = "DISABLED";
    FD1P3IX SLO__i16 (.D(SLO[14]), .SP(clk_enable_1114), .CD(GND_net), 
            .CK(clk), .Q(SLO[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i16.GSR = "DISABLED";
    FD1P3IX SLO__i19 (.D(SLO[17]), .SP(clk_enable_1114), .CD(GND_net), 
            .CK(clk), .Q(SLO[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i19.GSR = "DISABLED";
    FD1P3IX SLO__i13 (.D(SLO[11]), .SP(clk_enable_1114), .CD(GND_net), 
            .CK(clk), .Q(SLO[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i13.GSR = "DISABLED";
    FD1P3IX SLO__i17 (.D(SLO[15]), .SP(clk_enable_1114), .CD(GND_net), 
            .CK(clk), .Q(SLO[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i17.GSR = "DISABLED";
    FD1P3IX SLO__i20 (.D(SLO[18]), .SP(clk_enable_1114), .CD(GND_net), 
            .CK(clk), .Q(SLO[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i20.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_577 (.A(n27827), .B(\spi_data_out_r_39__N_5540[3] ), 
         .C(n3_adj_6704), .D(spi_data_out_r_39__N_5580), .Z(n27833)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_577.init = 16'hfefa;
    FD1P3IX SLO__i10 (.D(SLO[8]), .SP(clk_enable_1114), .CD(GND_net), 
            .CK(clk), .Q(SLO[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i10.GSR = "DISABLED";
    FD1P3IX SLO__i14 (.D(SLO[12]), .SP(clk_enable_1114), .CD(GND_net), 
            .CK(clk), .Q(SLO[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i14.GSR = "DISABLED";
    FD1P3IX SLO__i11 (.D(SLO[9]), .SP(clk_enable_1114), .CD(GND_net), 
            .CK(clk), .Q(SLO[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i11.GSR = "DISABLED";
    FD1P3IX SLO__i15 (.D(SLO[13]), .SP(clk_enable_1114), .CD(GND_net), 
            .CK(clk), .Q(SLO[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i15.GSR = "DISABLED";
    FD1P3IX SLO__i18 (.D(SLO[16]), .SP(clk_enable_1114), .CD(GND_net), 
            .CK(clk), .Q(SLO[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i18.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_578 (.A(\spi_data_out_r_39__N_4511[3] ), .B(n27823), 
         .C(n22_adj_6705), .D(spi_data_out_r_39__N_4551), .Z(n27831)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_578.init = 16'hfefc;
    LUT4 i1_4_lut_adj_579 (.A(\spi_data_out_r_39__N_1404[3] ), .B(\spi_data_out_r_39__N_1639[3] ), 
         .C(spi_data_out_r_39__N_1444), .D(spi_data_out_r_39__N_1679), .Z(n27817)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_579.init = 16'heca0;
    LUT4 i1_4_lut_adj_580 (.A(\spi_data_out_r_39__N_1874[3] ), .B(n27813), 
         .C(n8_adj_6706), .D(spi_data_out_r_39__N_1914), .Z(n27827)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_580.init = 16'hfefc;
    LUT4 Select_2911_i3_2_lut (.A(\spi_data_out_r_39__N_1169[3] ), .B(spi_data_out_r_39__N_1209), 
         .Z(n3_adj_6704)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2911_i3_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_581 (.A(\spi_data_out_r_39__N_2109[3] ), .B(\spi_data_out_r_39__N_934[3] ), 
         .C(spi_data_out_r_39__N_2149), .D(spi_data_out_r_39__N_974), .Z(n27813)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_581.init = 16'heca0;
    FD1P3IX SLO__i4 (.D(SLO[2]), .SP(clk_enable_1114), .CD(GND_net), .CK(clk), 
            .Q(SLO[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i4.GSR = "DISABLED";
    FD1P3IX SLO__i7 (.D(SLO[5]), .SP(clk_enable_1114), .CD(GND_net), .CK(clk), 
            .Q(SLO[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i7.GSR = "DISABLED";
    FD1P3IX SLO__i5 (.D(SLO[3]), .SP(clk_enable_1114), .CD(GND_net), .CK(clk), 
            .Q(SLO[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i5.GSR = "DISABLED";
    FD1P3IX SLO__i8 (.D(SLO[6]), .SP(clk_enable_1114), .CD(GND_net), .CK(clk), 
            .Q(SLO[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i8.GSR = "DISABLED";
    FD1P3IX SLO__i2 (.D(SLO[0]), .SP(clk_enable_1114), .CD(GND_net), .CK(clk), 
            .Q(SLO[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i2.GSR = "DISABLED";
    FD1P3IX SLO__i3 (.D(SLO[1]), .SP(clk_enable_1114), .CD(GND_net), .CK(clk), 
            .Q(SLO[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i3.GSR = "DISABLED";
    FD1P3IX SLO__i6 (.D(SLO[4]), .SP(clk_enable_1114), .CD(GND_net), .CK(clk), 
            .Q(SLO[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i6.GSR = "DISABLED";
    FD1P3IX SLO__i9 (.D(SLO[7]), .SP(clk_enable_1114), .CD(GND_net), .CK(clk), 
            .Q(SLO[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i9.GSR = "DISABLED";
    LUT4 Select_2911_i8_2_lut (.A(\spi_data_out_r_39__N_2344[3] ), .B(spi_data_out_r_39__N_2384), 
         .Z(n8_adj_6706)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2911_i8_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_582 (.A(\spi_data_out_r_39__N_5197[3] ), .B(\spi_data_out_r_39__N_4854[3] ), 
         .C(spi_data_out_r_39__N_5237), .D(spi_data_out_r_39__N_4894), .Z(n27823)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_582.init = 16'heca0;
    LUT4 Select_2911_i22_2_lut (.A(spi_data_out_r_39__N_5883[3]), .B(spi_data_out_r_39__N_5923), 
         .Z(n22_adj_6705)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_2911_i22_2_lut.init = 16'h8888;
    LUT4 SLO_buf_51__I_238_2_lut (.A(prev_MA_Temp), .B(MA_Temp), .Z(SLO_buf_51__N_6073)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[5:38])
    defparam SLO_buf_51__I_238_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_583 (.A(n27969), .B(n27977), .C(n27975), .D(n27961), 
         .Z(\spi_data_out_r[4] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_583.init = 16'hfffe;
    LUT4 i1_4_lut_adj_584 (.A(\spi_data_out_r_39__N_3825[4] ), .B(\spi_data_out_r_39__N_4168[4] ), 
         .C(spi_data_out_r_39__N_3865), .D(spi_data_out_r_39__N_4208), .Z(n27969)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_584.init = 16'heca0;
    FD1P3IX SLO__i1 (.D(pin_io_c_68), .SP(clk_enable_1114), .CD(GND_net), 
            .CK(clk), .Q(SLO[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=354, LSE_RLINE=397 */ ;   // c:/s_links/sources/slot_cards/stepper.v(129[8] 138[4])
    defparam SLO__i1.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_585 (.A(mode[0]), .B(mode[1]), .C(mode[2]), 
         .D(n30162), .Z(n26159)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_3_lut_4_lut_adj_585.init = 16'hfff7;
    LUT4 i24096_2_lut_3_lut (.A(mode[0]), .B(mode[1]), .C(mode[2]), .Z(ENC_O_N_6184)) /* synthesis lut_function=(!(A (B+(C))+!A (C))) */ ;
    defparam i24096_2_lut_3_lut.init = 16'h0707;
    LUT4 i24008_2_lut_rep_743 (.A(MA_Temp), .B(clk_1MHz), .Z(n30143)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i24008_2_lut_rep_743.init = 16'h7777;
    LUT4 i24172_2_lut_3_lut_4_lut (.A(MA_Temp), .B(clk_1MHz), .C(n30165), 
         .D(prev_MA), .Z(n12588)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i24172_2_lut_3_lut_4_lut.init = 16'h0007;
    LUT4 i1_2_lut_rep_665_3_lut (.A(MA_Temp), .B(clk_1MHz), .C(prev_MA), 
         .Z(n30065)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(118[13:34])
    defparam i1_2_lut_rep_665_3_lut.init = 16'hf8f8;
    
endmodule
//
// Verilog Description of module \uart_controller(DEV_ID=10,UART_ADDRESS_WIDTH=4) 
//

module \uart_controller(DEV_ID=10,UART_ADDRESS_WIDTH=4)  (uart_slot_en, clk, 
            clk_enable_320, n30185, \spi_data_r[0] , spi_cmd_r, n23978, 
            \spi_data_r[3] , \spi_data_r[2] , \spi_data_r[1] , \spi_addr_r[3] , 
            spi_data_valid_r, \spi_addr_r[0] , n26873, \spi_addr_r[1] , 
            n4, n23916) /* synthesis syn_module_defined=1 */ ;
    output [3:0]uart_slot_en;
    input clk;
    input clk_enable_320;
    input n30185;
    input \spi_data_r[0] ;
    input [15:0]spi_cmd_r;
    output n23978;
    input \spi_data_r[3] ;
    input \spi_data_r[2] ;
    input \spi_data_r[1] ;
    input \spi_addr_r[3] ;
    input spi_data_valid_r;
    input \spi_addr_r[0] ;
    output n26873;
    input \spi_addr_r[1] ;
    output n4;
    output n23916;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(70[18:21])
    
    wire n30171, n26867, n28436, n26855, n26851, n28500, n25509;
    
    FD1P3IX uart_slot_en_r__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_320), 
            .CD(n30185), .CK(clk), .Q(uart_slot_en[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=243, LSE_RLINE=254 */ ;   // c:/s_links/sources/uart_controller.v(57[8] 65[4])
    defparam uart_slot_en_r__i0.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(spi_cmd_r[9]), .B(spi_cmd_r[11]), .C(spi_cmd_r[14]), 
         .D(spi_cmd_r[13]), .Z(n23978)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut.init = 16'hfffe;
    FD1P3IX uart_slot_en_r__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_320), 
            .CD(n30185), .CK(clk), .Q(uart_slot_en[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=243, LSE_RLINE=254 */ ;   // c:/s_links/sources/uart_controller.v(57[8] 65[4])
    defparam uart_slot_en_r__i3.GSR = "DISABLED";
    FD1P3IX uart_slot_en_r__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_320), 
            .CD(n30185), .CK(clk), .Q(uart_slot_en[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=243, LSE_RLINE=254 */ ;   // c:/s_links/sources/uart_controller.v(57[8] 65[4])
    defparam uart_slot_en_r__i2.GSR = "DISABLED";
    FD1P3IX uart_slot_en_r__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_320), 
            .CD(n30185), .CK(clk), .Q(uart_slot_en[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=243, LSE_RLINE=254 */ ;   // c:/s_links/sources/uart_controller.v(57[8] 65[4])
    defparam uart_slot_en_r__i1.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_771 (.A(\spi_addr_r[3] ), .B(spi_data_valid_r), .Z(n30171)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_771.init = 16'h8888;
    LUT4 i1_4_lut_adj_304 (.A(\spi_addr_r[0] ), .B(n23978), .C(n26867), 
         .D(spi_cmd_r[3]), .Z(n26873)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_304.init = 16'h0010;
    LUT4 i1_4_lut_adj_305 (.A(n28436), .B(spi_cmd_r[7]), .C(n26855), .D(spi_cmd_r[8]), 
         .Z(n26867)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_305.init = 16'h0010;
    LUT4 i23734_4_lut (.A(spi_cmd_r[12]), .B(spi_cmd_r[6]), .C(spi_cmd_r[10]), 
         .D(spi_cmd_r[15]), .Z(n28436)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23734_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_306 (.A(spi_cmd_r[2]), .B(n26851), .C(n30171), .D(spi_cmd_r[4]), 
         .Z(n26855)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_306.init = 16'h8000;
    LUT4 i1_2_lut (.A(spi_cmd_r[1]), .B(spi_cmd_r[5]), .Z(n26851)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_307 (.A(\spi_addr_r[1] ), .B(spi_cmd_r[0]), .Z(n4)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_307.init = 16'h2222;
    LUT4 i1_4_lut_adj_308 (.A(n28500), .B(n23978), .C(n25509), .D(spi_cmd_r[7]), 
         .Z(n23916)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_4_lut_adj_308.init = 16'h0010;
    LUT4 i23798_4_lut (.A(spi_cmd_r[12]), .B(spi_cmd_r[10]), .C(spi_cmd_r[6]), 
         .D(spi_cmd_r[8]), .Z(n28500)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i23798_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_309 (.A(spi_cmd_r[15]), .B(spi_data_valid_r), .Z(n25509)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_309.init = 16'h4444;
    
endmodule
