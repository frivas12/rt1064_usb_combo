// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.12.0.240.2
// Netlist written on Mon Apr 11 16:49:49 2022
//
// Verilog Description of module mcm_top
//

module mcm_top (clk_in, resetn, led_sw, cs, intrpt_out, FLASH_CS, 
            MAX3421_CS, CS_READY, spi_clk, spi_mosi, spi_miso, spi_scsn, 
            UC_TXD0, UC_RXD0, pin_io, C_1, C_2, C_3, C_4, C_5, 
            C_6, C_7, C_8) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(9[8:15])
    input clk_in;   // c:/s_links/sources/mcm_top.v(16[27:33])
    input resetn;   // c:/s_links/sources/mcm_top.v(17[27:33])
    output led_sw;   // c:/s_links/sources/mcm_top.v(18[24:30])
    input [4:0]cs;   // c:/s_links/sources/mcm_top.v(19[37:39])
    output [6:0]intrpt_out;   // c:/s_links/sources/mcm_top.v(20[36:46])
    output FLASH_CS;   // c:/s_links/sources/mcm_top.v(21[24:32])
    output MAX3421_CS;   // c:/s_links/sources/mcm_top.v(22[24:34])
    input CS_READY;   // c:/s_links/sources/mcm_top.v(23[24:32])
    input spi_clk /* synthesis black_box_pad_pin=1 */ ;   // c:/s_links/sources/mcm_top.v(26[27:34])
    input spi_mosi /* synthesis black_box_pad_pin=1 */ ;   // c:/s_links/sources/mcm_top.v(27[27:35])
    output spi_miso /* synthesis black_box_pad_pin=1 */ ;   // c:/s_links/sources/mcm_top.v(28[27:35])
    input spi_scsn;   // c:/s_links/sources/mcm_top.v(29[27:35])
    input UC_TXD0;   // c:/s_links/sources/mcm_top.v(32[27:34])
    output UC_RXD0;   // c:/s_links/sources/mcm_top.v(33[27:34])
    inout [69:0]pin_io;   // c:/s_links/sources/mcm_top.v(36[51:57])
    output C_1 /* synthesis .original_dir=IN_OUT */ ;   // c:/s_links/sources/mcm_top.v(39[24:27])
    output C_2 /* synthesis .original_dir=IN_OUT */ ;   // c:/s_links/sources/mcm_top.v(40[24:27])
    output C_3 /* synthesis .original_dir=IN_OUT */ ;   // c:/s_links/sources/mcm_top.v(41[24:27])
    output C_4 /* synthesis .original_dir=IN_OUT */ ;   // c:/s_links/sources/mcm_top.v(42[24:27])
    output C_5 /* synthesis .original_dir=IN_OUT */ ;   // c:/s_links/sources/mcm_top.v(43[24:27])
    inout C_6;   // c:/s_links/sources/mcm_top.v(44[24:27])
    output C_7 /* synthesis .original_dir=IN_OUT */ ;   // c:/s_links/sources/mcm_top.v(45[24:27])
    input C_8 /* synthesis .original_dir=IN_OUT */ ;   // c:/s_links/sources/mcm_top.v(46[24:27])
    
    wire clk_in_c /* synthesis is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(16[27:33])
    wire CS_READY_c /* synthesis is_clock=1, SET_AS_NETWORK=CS_READY_c */ ;   // c:/s_links/sources/mcm_top.v(23[24:32])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire [20:0]pin_intrpt /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[20] */ ;   // c:/s_links/sources/mcm_top.v(102[46:56])
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire mode_2_derived_32 /* synthesis is_clock=1, SET_AS_NETWORK=\stepper_ins[0].u_stepper/mode[2]_derived_32 */ ;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    wire mode_2_derived_32_adj_8013 /* synthesis is_clock=1, SET_AS_NETWORK=\stepper_ins[2].u_stepper/mode[2]_derived_32 */ ;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    wire mode_2_derived_32_adj_8049 /* synthesis is_clock=1, SET_AS_NETWORK=\stepper_ins[5].u_stepper/mode[2]_derived_32 */ ;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    wire spi_clk_i /* synthesis is_clock=1 */ ;   // c:/s_links/sources/config_mcm/ip/spi_slave_efb.v(34[10:19])
    
    wire GND_net, resetn_c, led_sw_c, cs_c_4, cs_c_3, cs_c_2, cs_c_1, 
        cs_c_0, intrpt_out_c_6, intrpt_out_c_5, intrpt_out_c_4, intrpt_out_c_3, 
        intrpt_out_c_2, intrpt_out_c_1, intrpt_out_c_0, FLASH_CS_c, 
        MAX3421_CS_c, spi_scsn_c, C_5_c_c, n19, n15, n13, n11, 
        n8, n4, n7, C_1_c_0, C_2_c_1, C_3_c_2, C_4_c_3, C_8_c;
    wire [15:0]spi_cmd_r;   // c:/s_links/sources/mcm_top.v(83[27:36])
    wire [7:0]spi_addr_r;   // c:/s_links/sources/mcm_top.v(84[28:38])
    wire [39:0]spi_data_r;   // c:/s_links/sources/mcm_top.v(85[22:32])
    
    wire spi_data_valid_r;
    wire [15:0]spi_cmd;   // c:/s_links/sources/mcm_top.v(88[27:34])
    wire [7:0]spi_addr;   // c:/s_links/sources/mcm_top.v(89[28:36])
    wire [39:0]spi_data_out_r;   // c:/s_links/sources/mcm_top.v(90[22:36])
    wire [13:0]cs_decoded;   // c:/s_links/sources/mcm_top.v(93[43:53])
    wire [6:0]quad_a;   // c:/s_links/sources/mcm_top.v(98[31:37])
    wire [6:0]quad_b;   // c:/s_links/sources/mcm_top.v(99[31:37])
    
    wire EM_STOP, n27286, spi_cmd_valid, spi_addr_valid, spi_data_valid, 
        spi_sdo_valid_N_297, n29075, n65, spi_sdo_valid_N_296, n26969, 
        n6, clk_enable_288, clk_1MHz_enable_367, n29091, n26525, n29256, 
        n2;
    wire [39:0]spi_data_out_r_39__N_770;
    
    wire spi_data_out_r_39__N_810;
    wire [1:0]quad_homing;   // c:/s_links/sources/quad_decoder.v(41[19:30])
    
    wire quad_set_valid, quad_set_complete, n27058;
    wire [39:0]spi_data_out_r_39__N_934;
    
    wire spi_data_out_r_39__N_1162, spi_data_out_r_39__N_974, n29255, 
        clk_enable_400, n29254, clk_enable_505, n26579, n29251;
    wire [1:0]quad_homing_adj_8225;   // c:/s_links/sources/quad_decoder.v(41[19:30])
    
    wire quad_set_complete_adj_7619;
    wire [31:0]quad_count_adj_8226;   // c:/s_links/sources/quad_decoder.v(45[29:39])
    wire [31:0]quad_buffer_adj_8227;   // c:/s_links/sources/quad_decoder.v(46[29:40])
    
    wire clk_1MHz_enable_40, n26951, clk_enable_526;
    wire [39:0]spi_data_out_r_39__N_1313;
    wire [39:0]spi_data_out_r_39__N_1168;
    
    wire spi_data_out_r_39__N_1396, spi_data_out_r_39__N_1208, n29247, 
        n26569, n2_adj_7620;
    wire [1:0]quad_homing_adj_8284;   // c:/s_links/sources/quad_decoder.v(41[19:30])
    
    wire quad_set_complete_adj_7623;
    wire [31:0]quad_count_adj_8285;   // c:/s_links/sources/quad_decoder.v(45[29:39])
    wire [31:0]quad_buffer_adj_8286;   // c:/s_links/sources/quad_decoder.v(46[29:40])
    wire [39:0]spi_data_out_r_39__N_1547;
    
    wire n47, n26565;
    wire [39:0]spi_data_out_r_39__N_1402;
    
    wire spi_data_out_r_39__N_1442, n29089, n13265, n22, n26561;
    wire [1:0]quad_homing_adj_8343;   // c:/s_links/sources/quad_decoder.v(41[19:30])
    
    wire quad_set_complete_adj_7689;
    wire [31:0]quad_count_adj_8344;   // c:/s_links/sources/quad_decoder.v(45[29:39])
    wire [31:0]quad_buffer_adj_8345;   // c:/s_links/sources/quad_decoder.v(46[29:40])
    
    wire n19084, n24, n29239;
    wire [39:0]spi_data_out_r_39__N_1781;
    wire [39:0]spi_data_out_r_39__N_1636;
    
    wire spi_data_out_r_39__N_1676, n29237, n32, n22_adj_7754, n19233, 
        n29233, n26549, n27338, n29336, n25411, n3, n29225;
    wire [1:0]quad_homing_adj_8402;   // c:/s_links/sources/quad_decoder.v(41[19:30])
    
    wire quad_set_complete_adj_7757;
    wire [31:0]quad_count_adj_8403;   // c:/s_links/sources/quad_decoder.v(45[29:39])
    wire [31:0]quad_buffer_adj_8404;   // c:/s_links/sources/quad_decoder.v(46[29:40])
    
    wire clk_enable_359, clk_1MHz_enable_66, n29224;
    wire [39:0]spi_data_out_r_39__N_2015;
    wire [39:0]spi_data_out_r_39__N_1870;
    
    wire spi_data_out_r_39__N_2098, spi_data_out_r_39__N_1910, clk_enable_206, 
        clk_enable_190, n29220;
    wire [1:0]quad_homing_adj_8461;   // c:/s_links/sources/quad_decoder.v(41[19:30])
    
    wire quad_set_valid_adj_7824, quad_set_complete_adj_7825;
    wire [31:0]quad_count_adj_8462;   // c:/s_links/sources/quad_decoder.v(45[29:39])
    wire [31:0]quad_buffer_adj_8463;   // c:/s_links/sources/quad_decoder.v(46[29:40])
    
    wire n26, n26938, n29217, n29216, n31, n26521;
    wire [39:0]spi_data_out_r_39__N_2249;
    wire [39:0]spi_data_out_r_39__N_2104;
    
    wire spi_data_out_r_39__N_2332, spi_data_out_r_39__N_2144, clk_enable_188, 
        clk_enable_174, clk_enable_177, clk_enable_183, clk_enable_185, 
        clk_enable_187, clk_enable_192, clk_enable_194, clk_enable_193, 
        clk_enable_204, clk_enable_200, clk_enable_32, clk_enable_172, 
        clk_enable_169, clk_enable_171, clk_enable_176, clk_enable_179, 
        clk_enable_189, clk_enable_191, clk_enable_182, clk_enable_166, 
        clk_enable_201, clk_enable_202, clk_enable_197, clk_enable_167, 
        clk_enable_170, clk_enable_175, clk_enable_178, n29214, n13_adj_7890, 
        quad_set_complete_adj_7891;
    wire [31:0]quad_count_adj_8521;   // c:/s_links/sources/quad_decoder.v(45[29:39])
    wire [31:0]quad_buffer_adj_8522;   // c:/s_links/sources/quad_decoder.v(46[29:40])
    
    wire n27283, n13052, n29213, n29212, n29211;
    wire [39:0]spi_data_out_r_39__N_2483;
    wire [39:0]spi_data_out_r_39__N_2338;
    
    wire spi_data_out_r_39__N_2566, spi_data_out_r_39__N_2378, clk_enable_86, 
        n27480, clk_1MHz_enable_182, clk_enable_180, clk_enable_181, 
        clk_enable_184, clk_enable_186, n29210, clk_enable_20, n29207, 
        n27471, n26972, n8826, clear_intrpt, clear_intrpt_N_2639, 
        n26529, n29205, n5;
    wire [39:0]spi_data_out_r_39__N_2572;
    
    wire intrpt_out_N_2635, n26523, clear_intrpt_adj_7956, clear_intrpt_N_2710, 
        n2_adj_7957;
    wire [39:0]spi_data_out_r_39__N_2643;
    
    wire intrpt_out_N_2706, clear_intrpt_adj_7958, clear_intrpt_N_2781;
    wire [39:0]spi_data_out_r_39__N_2714;
    
    wire intrpt_out_N_2777, clear_intrpt_adj_7959, clear_intrpt_N_2852, 
        n29204, n29203;
    wire [39:0]spi_data_out_r_39__N_2785;
    
    wire intrpt_out_N_2848, clear_intrpt_adj_7960, clear_intrpt_N_2923, 
        n29202;
    wire [39:0]spi_data_out_r_39__N_2856;
    
    wire intrpt_out_N_2919, clear_intrpt_adj_7961, n29201, clear_intrpt_N_2994, 
        n29200;
    wire [39:0]spi_data_out_r_39__N_2927;
    
    wire intrpt_out_N_2990, clear_intrpt_adj_7962, clear_intrpt_N_3065, 
        n29199;
    wire [39:0]spi_data_out_r_39__N_2998;
    
    wire intrpt_out_N_3061, n29198, clk_enable_164, clk_enable_271, 
        clk_1MHz_enable_24, n29196, n29195, n29194, clk_enable_30, 
        clk_1MHz_enable_91, n29193, n27657, n27465, n27477, n27301, 
        n29191, n29190, n29189, n27590, n27234, clk_enable_402, 
        clk_1MHz_enable_55, clk_enable_76, clk_enable_499, n29185, clk_enable_131, 
        clk_enable_28, n3_adj_7963, clk_enable_162, clk_enable_77;
    wire [2:0]n29780;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    wire reset_r, digital_output_r, n27189, n26533, n2_adj_7964, n12716, 
        n29182;
    wire [39:0]spi_data_out_r_39__N_3818;
    
    wire spi_data_out_r_39__N_3858, n2_adj_7965;
    wire [2:0]n29781;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    wire reset_r_adj_7969, digital_output_r_adj_7970;
    wire [51:0]SLO_buf_adj_8796;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire OW_ID_N_4464, OW_ID_N_4462, n26535, n2_adj_7971, n9633, reset_r_N_4474;
    wire [39:0]spi_data_out_r_39__N_4419;
    wire [39:0]spi_data_out_r_39__N_4157;
    
    wire spi_data_out_r_39__N_4490, spi_data_out_r_39__N_4197;
    wire [2:0]n29782;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    wire reset_r_adj_7975, digital_output_r_adj_7976, clk_enable_398, 
        n2_adj_7977, n29326, n29178, n18550, reset_r_N_4813;
    wire [39:0]spi_data_out_r_39__N_4496;
    
    wire spi_data_out_r_39__N_4536;
    wire [2:0]n29783;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    wire reset_r_adj_7981, digital_output_r_adj_7982, NSL, clk_enable_199;
    wire [51:0]SLO_buf_adj_8858;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire clk_enable_434, n19401, n29174, n27240, n13615, n19391, 
        n19381, clk_enable_340;
    wire [39:0]spi_data_out_r_39__N_5097;
    wire [39:0]spi_data_out_r_39__N_4835;
    
    wire spi_data_out_r_39__N_4875, n13511;
    wire [2:0]n29784;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    wire reset_r_adj_8017, digital_output_r_adj_8018;
    wire [51:0]SLO_buf_adj_8889;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire OW_ID_N_5482, n29087, n26531, n13413, n19371;
    wire [39:0]spi_data_out_r_39__N_5436;
    wire [39:0]spi_data_out_r_39__N_5174;
    
    wire spi_data_out_r_39__N_5507, spi_data_out_r_39__N_5214;
    wire [2:0]n29785;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    wire reset_r_adj_8053, digital_output_r_adj_8054, n13489, n29169;
    wire [51:0]SLO_buf_adj_8920;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire n19361, n28813, n28811, n13506, n19351, n31_adj_8085;
    wire [39:0]spi_data_out_r_39__N_5775;
    wire [39:0]spi_data_out_r_39__N_5513;
    
    wire spi_data_out_r_39__N_5553;
    wire [2:0]n29786;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    wire reset_r_adj_8089, digital_output_r_adj_8090;
    wire [51:0]SLO_buf_adj_8951;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire n19337, n6_adj_8121;
    wire [39:0]spi_data_out_r_39__N_6114;
    wire [39:0]spi_data_out_r_39__N_5852;
    
    wire spi_data_out_r_39__N_5892, VCC_net, mode, n13074, mode_adj_8122, 
        mode_adj_8123, mode_adj_8124, mode_adj_8125, clk_enable_198, 
        mode_adj_8126, mode_adj_8127, n29162, n29161, mode_adj_8128, 
        mode_adj_8129, n29160, n27483, n29158, mode_adj_8130, n27618, 
        mode_adj_8131, n29157, mode_adj_8132, mode_adj_8133, mode_adj_8134, 
        mode_adj_8135, n5_adj_8136, n29153, mode_adj_8137, n29070, 
        n1, mode_adj_8138, mode_adj_8139, mode_adj_8140, mode_adj_8141, 
        mode_adj_8142, mode_adj_8143, clk_enable_173, tx_N_6443, n26963, 
        mode_adj_8144, mode_adj_8145, clk_enable_269, mode_adj_8146, 
        mode_adj_8147, n29150, mode_adj_8148, n29149, mode_adj_8149, 
        mode_adj_8150, spi_mosi_oe, spi_mosi_o, spi_miso_oe, spi_miso_o, 
        spi_clk_oe, spi_clk_o, spi_mosi_i, spi_miso_i, mem_rdata_update_N_729, 
        clk_enable_435, clk_enable_467, clk_enable_286, n29144, n27225, 
        clk_enable_433, clk_enable_436, clk_enable_509, n29141, clk_enable_303, 
        n12714, clk_enable_524, n25293, n13_adj_8151, n5647, n27259, 
        n27, n29757, n65_adj_8152, n31_adj_8153, n21446, n29085, 
        clk_enable_503, n29134, n29132, n29084, n66, n29130, n20819, 
        n95, n29127, n29126, clk_enable_501, n14, n26928, n27632, 
        n26948, clk_1MHz_enable_171, n29124, n27186, n27636, n29123, 
        n29083, n29762, clk_enable_502, n29122, n29761, n79, clk_enable_307, 
        clk_enable_506, n29120, clk_enable_519, clk_1MHz_enable_340, 
        clk_enable_520, n29118, n29117, n108, n25382, n29317, n29315, 
        n29313, n29311, n29310, n29115, n29309, n29307, n29306, 
        n29305, n29303, n29301, n29114, n29300, n27285, clk_enable_518, 
        n29299, n26965, n29110, n29295, n1_adj_8154, n2_adj_8155, 
        n8633, n29293, n1_adj_8156, n1_adj_8157, n8651, n8652, n1_adj_8158, 
        n2_adj_8159, n8661, n29108, n29106, n1_adj_8160, n1_adj_8161, 
        n8679, n8680, n1_adj_8162, n2_adj_8163, n8689, n27256, clk_enable_306, 
        n29105, n1_adj_8164, n1_adj_8165, n29104, n8716, n8717, 
        n2_adj_8166, n8720, n29102, n1_adj_8167, pin_io_out_69, n1_adj_8168, 
        n8739, n8740, n1_adj_8169, n2_adj_8170, n8749, n1_adj_8171, 
        n1_adj_8172, n8767, n8768, n1_adj_8173, n2_adj_8174, n8777, 
        n29288, n1_adj_8175, n1_adj_8176, n8795, n8796, n1_adj_8177, 
        n29287, n2_adj_8178, n8805, clk_enable_342, n29101, n1_adj_8179, 
        n29100, n8823, n8824, pin_io_out_68, pin_io_out_66, pin_io_out_65, 
        pin_io_out_64, n29286, pin_io_out_63, n8836, pin_io_out_62, 
        n29099, pin_io_out_59, n8840, pin_io_out_58, pin_io_out_56, 
        pin_io_out_55, pin_io_out_54, pin_io_out_53, n8850, pin_io_out_52, 
        n29098, pin_io_out_49, n8854, pin_io_out_48, pin_io_out_46, 
        pin_io_out_45, pin_io_out_44, pin_io_out_43, n8864, pin_io_out_42, 
        pin_io_out_40, pin_io_out_39, n8870, pin_io_out_38, pin_io_out_36, 
        pin_io_out_35, pin_io_out_34, n29285, pin_io_out_33, n8880, 
        pin_io_out_32, pin_io_out_29, n8884, pin_io_out_28, pin_io_out_26, 
        pin_io_out_25, pin_io_out_24, pin_io_out_23, n8894, pin_io_out_22, 
        pin_io_out_19, n8898, pin_io_out_18, pin_io_out_16, pin_io_out_15, 
        pin_io_out_14, pin_io_out_13, n8908, pin_io_out_12, pin_io_out_9, 
        pin_io_out_8, pin_io_out_6, pin_io_out_5, pin_io_out_4, pin_io_out_3, 
        n8922, pin_io_out_2, UC_RXD0_c, n29284, n29282, n2_adj_8180, 
        n3_adj_8181, n4_adj_8182, n11_adj_8183, n15_adj_8184, n17, 
        n29097, n29096, n20, n21, n29082, n29080, n29079, n29078, 
        n29077, n29076, n29094, n29267, clk_enable_521, n29093, 
        n29092, n26933, n29260;
    
    VHI i2 (.Z(VCC_net));
    BB BBspi_mosi (.I(spi_mosi_o), .T(spi_mosi_oe), .B(spi_mosi), .O(spi_mosi_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=15, LSE_LLINE=162, LSE_RLINE=176 */ ;   // c:/s_links/sources/config_mcm/ip/spi_slave_efb.v(39[8:82])
    OSCH OSCH_inst (.STDBY(GND_net), .OSC(clk)) /* synthesis syn_instantiated=1 */ ;
    defparam OSCH_inst.NOM_FREQ = "38.00";
    BB BBspi_miso (.I(spi_miso_o), .T(spi_miso_oe), .B(spi_miso), .O(spi_miso_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=15, LSE_LLINE=162, LSE_RLINE=176 */ ;   // c:/s_links/sources/config_mcm/ip/spi_slave_efb.v(41[8:82])
    BB BBspi_clk (.I(spi_clk_o), .T(spi_clk_oe), .B(spi_clk), .O(spi_clk_i)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=15, LSE_LLINE=162, LSE_RLINE=176 */ ;   // c:/s_links/sources/config_mcm/ip/spi_slave_efb.v(43[8:77])
    IB C_8_pad (.I(C_8), .O(C_8_c));   // c:/s_links/sources/mcm_top.v(46[24:27])
    IB C_5_c_pad (.I(UC_TXD0), .O(C_5_c_c));   // c:/s_links/sources/mcm_top.v(32[27:34])
    IB spi_scsn_pad (.I(spi_scsn), .O(spi_scsn_c));   // c:/s_links/sources/mcm_top.v(29[27:35])
    IB CS_READY_pad (.I(CS_READY), .O(CS_READY_c));   // c:/s_links/sources/mcm_top.v(23[24:32])
    IB cs_pad_0 (.I(cs[0]), .O(cs_c_0));   // c:/s_links/sources/mcm_top.v(19[37:39])
    IB cs_pad_1 (.I(cs[1]), .O(cs_c_1));   // c:/s_links/sources/mcm_top.v(19[37:39])
    IB cs_pad_2 (.I(cs[2]), .O(cs_c_2));   // c:/s_links/sources/mcm_top.v(19[37:39])
    IB cs_pad_3 (.I(cs[3]), .O(cs_c_3));   // c:/s_links/sources/mcm_top.v(19[37:39])
    IB cs_pad_4 (.I(cs[4]), .O(cs_c_4));   // c:/s_links/sources/mcm_top.v(19[37:39])
    IB resetn_pad (.I(resetn), .O(resetn_c));   // c:/s_links/sources/mcm_top.v(17[27:33])
    IB clk_in_pad (.I(clk_in), .O(clk_in_c));   // c:/s_links/sources/mcm_top.v(16[27:33])
    OBZ C_7_pad (.I(C_5_c_c), .T(tx_N_6443), .O(C_7));   // c:/s_links/sources/slot_cards/peizo_elliptec.v(30[8:10])
    OB C_5_pad (.I(C_5_c_c), .O(C_5));   // c:/s_links/sources/mcm_top.v(43[24:27])
    OB C_4_pad (.I(C_4_c_3), .O(C_4));   // c:/s_links/sources/mcm_top.v(42[24:27])
    OB C_3_pad (.I(C_3_c_2), .O(C_3));   // c:/s_links/sources/mcm_top.v(41[24:27])
    OB C_2_pad (.I(C_2_c_1), .O(C_2));   // c:/s_links/sources/mcm_top.v(40[24:27])
    OB C_1_pad (.I(C_1_c_0), .O(C_1));   // c:/s_links/sources/mcm_top.v(39[24:27])
    OBZ pin_io_pad_0 (.I(n8824), .T(n8823), .O(pin_io[0]));
    OBZ pin_io_pad_1 (.I(n1_adj_8179), .T(n29260), .O(pin_io[1]));
    OBZ pin_io_pad_7 (.I(n1_adj_8177), .T(n29185), .O(pin_io[7]));
    OBZ pin_io_pad_10 (.I(n8796), .T(n8795), .O(pin_io[10]));
    OBZ pin_io_pad_11 (.I(n1_adj_8175), .T(n29237), .O(pin_io[11]));
    OBZ pin_io_pad_17 (.I(n1_adj_8173), .T(n29217), .O(pin_io[17]));
    OBZ pin_io_pad_20 (.I(n8768), .T(n8767), .O(pin_io[20]));
    OBZ pin_io_pad_21 (.I(n1_adj_8171), .T(n29233), .O(pin_io[21]));
    OBZ pin_io_pad_27 (.I(n1_adj_8169), .T(n29295), .O(pin_io[27]));
    OBZ pin_io_pad_30 (.I(n8740), .T(n8739), .O(pin_io[30]));
    OBZ pin_io_pad_31 (.I(n1_adj_8167), .T(n29225), .O(pin_io[31]));
    OBZ pin_io_pad_37 (.I(n8717), .T(n8716), .O(pin_io[37]));
    OBZ pin_io_pad_41 (.I(n1_adj_8164), .T(n29224), .O(pin_io[41]));
    OBZ pin_io_pad_47 (.I(n1_adj_8162), .T(n29207), .O(pin_io[47]));
    OBZ pin_io_pad_50 (.I(n8680), .T(n8679), .O(pin_io[50]));
    OBZ pin_io_pad_51 (.I(n1_adj_8160), .T(n29220), .O(pin_io[51]));
    OBZ pin_io_pad_57 (.I(n1_adj_8158), .T(n29210), .O(pin_io[57]));
    OBZ pin_io_pad_60 (.I(n8652), .T(n8651), .O(pin_io[60]));
    OBZ pin_io_pad_61 (.I(n1_adj_8156), .T(n29267), .O(pin_io[61]));
    OBZ pin_io_pad_67 (.I(n1_adj_8154), .T(n29195), .O(pin_io[67]));
    OB UC_RXD0_pad (.I(UC_RXD0_c), .O(UC_RXD0));   // c:/s_links/sources/mcm_top.v(33[27:34])
    OB MAX3421_CS_pad (.I(MAX3421_CS_c), .O(MAX3421_CS));   // c:/s_links/sources/mcm_top.v(22[24:34])
    OB FLASH_CS_pad (.I(FLASH_CS_c), .O(FLASH_CS));   // c:/s_links/sources/mcm_top.v(21[24:32])
    OB intrpt_out_pad_0 (.I(intrpt_out_c_0), .O(intrpt_out[0]));   // c:/s_links/sources/mcm_top.v(20[36:46])
    OB intrpt_out_pad_1 (.I(intrpt_out_c_1), .O(intrpt_out[1]));   // c:/s_links/sources/mcm_top.v(20[36:46])
    OB intrpt_out_pad_2 (.I(intrpt_out_c_2), .O(intrpt_out[2]));   // c:/s_links/sources/mcm_top.v(20[36:46])
    OB intrpt_out_pad_3 (.I(intrpt_out_c_3), .O(intrpt_out[3]));   // c:/s_links/sources/mcm_top.v(20[36:46])
    OB intrpt_out_pad_4 (.I(intrpt_out_c_4), .O(intrpt_out[4]));   // c:/s_links/sources/mcm_top.v(20[36:46])
    OB intrpt_out_pad_5 (.I(intrpt_out_c_5), .O(intrpt_out[5]));   // c:/s_links/sources/mcm_top.v(20[36:46])
    OB intrpt_out_pad_6 (.I(intrpt_out_c_6), .O(intrpt_out[6]));   // c:/s_links/sources/mcm_top.v(20[36:46])
    OB led_sw_pad (.I(led_sw_c), .O(led_sw));   // c:/s_links/sources/mcm_top.v(18[24:30])
    BB UC_RXD0_pad_4167 (.I(n25382), .T(n26951), .B(C_6), .O(UC_RXD0_c));
    BB pin_io_pad_2 (.I(GND_net), .T(VCC_net), .B(pin_io[2]), .O(pin_io_out_2));   // c:/s_links/sources/slot_cards/shutter_4.v(68[8:14])
    BB pin_io_pad_3 (.I(n2_adj_8178), .T(n8922), .B(pin_io[3]), .O(pin_io_out_3));
    BB pin_io_pad_4 (.I(GND_net), .T(VCC_net), .B(pin_io[4]), .O(pin_io_out_4));   // c:/s_links/sources/slot_cards/shutter_4.v(70[8:14])
    BB pin_io_pad_5 (.I(n26535), .T(n26561), .B(pin_io[5]), .O(pin_io_out_5));
    BB pin_io_pad_6 (.I(n2_adj_7977), .T(n8805), .B(pin_io[6]), .O(pin_io_out_6));
    BB pin_io_pad_8 (.I(GND_net), .T(VCC_net), .B(pin_io[8]), .O(pin_io_out_8));   // c:/s_links/sources/slot_cards/shutter_4.v(73[8:14])
    BB pin_io_pad_9 (.I(n1_adj_8176), .T(n3_adj_7963), .B(pin_io[9]), 
       .O(pin_io_out_9));
    BB pin_io_pad_12 (.I(GND_net), .T(VCC_net), .B(pin_io[12]), .O(pin_io_out_12));   // c:/s_links/sources/slot_cards/shutter_4.v(68[8:14])
    BB pin_io_pad_13 (.I(n2_adj_8174), .T(n8908), .B(pin_io[13]), .O(pin_io_out_13));
    BB pin_io_pad_14 (.I(GND_net), .T(VCC_net), .B(pin_io[14]), .O(pin_io_out_14));   // c:/s_links/sources/slot_cards/shutter_4.v(70[8:14])
    BB pin_io_pad_15 (.I(n26533), .T(n13615), .B(pin_io[15]), .O(pin_io_out_15));
    BB pin_io_pad_16 (.I(n2_adj_7971), .T(n8777), .B(pin_io[16]), .O(pin_io_out_16));
    BB pin_io_pad_18 (.I(GND_net), .T(VCC_net), .B(pin_io[18]), .O(pin_io_out_18));   // c:/s_links/sources/slot_cards/shutter_4.v(73[8:14])
    BB pin_io_pad_19 (.I(n1_adj_8172), .T(n8898), .B(pin_io[19]), .O(pin_io_out_19));
    BB pin_io_pad_22 (.I(GND_net), .T(VCC_net), .B(pin_io[22]), .O(pin_io_out_22));   // c:/s_links/sources/slot_cards/shutter_4.v(68[8:14])
    BB pin_io_pad_23 (.I(n2_adj_8170), .T(n8894), .B(pin_io[23]), .O(pin_io_out_23));
    BB pin_io_pad_24 (.I(GND_net), .T(VCC_net), .B(pin_io[24]), .O(pin_io_out_24));   // c:/s_links/sources/slot_cards/shutter_4.v(70[8:14])
    BB pin_io_pad_25 (.I(n26531), .T(n26549), .B(pin_io[25]), .O(pin_io_out_25));
    BB pin_io_pad_26 (.I(n2_adj_7964), .T(n8749), .B(pin_io[26]), .O(pin_io_out_26));
    BB pin_io_pad_28 (.I(GND_net), .T(VCC_net), .B(pin_io[28]), .O(pin_io_out_28));   // c:/s_links/sources/slot_cards/shutter_4.v(73[8:14])
    BB pin_io_pad_29 (.I(n1_adj_8168), .T(n8884), .B(pin_io[29]), .O(pin_io_out_29));
    BB pin_io_pad_32 (.I(GND_net), .T(VCC_net), .B(pin_io[32]), .O(pin_io_out_32));   // c:/s_links/sources/slot_cards/shutter_4.v(68[8:14])
    BB pin_io_pad_33 (.I(n2_adj_8166), .T(n8880), .B(pin_io[33]), .O(pin_io_out_33));
    BB pin_io_pad_34 (.I(GND_net), .T(VCC_net), .B(pin_io[34]), .O(pin_io_out_34));   // c:/s_links/sources/slot_cards/shutter_4.v(70[8:14])
    BB pin_io_pad_35 (.I(n26529), .T(n26565), .B(pin_io[35]), .O(pin_io_out_35));
    BB pin_io_pad_36 (.I(n2_adj_7957), .T(n8720), .B(pin_io[36]), .O(pin_io_out_36));
    BB pin_io_pad_38 (.I(GND_net), .T(VCC_net), .B(pin_io[38]), .O(pin_io_out_38));   // c:/s_links/sources/slot_cards/shutter_4.v(73[8:14])
    BB pin_io_pad_39 (.I(n1_adj_8165), .T(n8870), .B(pin_io[39]), .O(pin_io_out_39));
    BB pin_io_pad_40 (.I(n26965), .T(n25411), .B(pin_io[40]), .O(pin_io_out_40));
    BB pin_io_pad_42 (.I(GND_net), .T(VCC_net), .B(pin_io[42]), .O(pin_io_out_42));   // c:/s_links/sources/slot_cards/shutter_4.v(68[8:14])
    BB pin_io_pad_43 (.I(n2_adj_8163), .T(n8864), .B(pin_io[43]), .O(pin_io_out_43));
    BB pin_io_pad_44 (.I(GND_net), .T(VCC_net), .B(pin_io[44]), .O(pin_io_out_44));   // c:/s_links/sources/slot_cards/shutter_4.v(70[8:14])
    BB pin_io_pad_45 (.I(n26525), .T(n26569), .B(pin_io[45]), .O(pin_io_out_45));
    BB pin_io_pad_46 (.I(n2), .T(n8689), .B(pin_io[46]), .O(pin_io_out_46));
    BB pin_io_pad_48 (.I(GND_net), .T(VCC_net), .B(pin_io[48]), .O(pin_io_out_48));   // c:/s_links/sources/slot_cards/shutter_4.v(73[8:14])
    BB pin_io_pad_49 (.I(n1_adj_8161), .T(n8854), .B(pin_io[49]), .O(pin_io_out_49));
    BB pin_io_pad_52 (.I(GND_net), .T(VCC_net), .B(pin_io[52]), .O(pin_io_out_52));   // c:/s_links/sources/slot_cards/shutter_4.v(68[8:14])
    BB pin_io_pad_53 (.I(n2_adj_8159), .T(n8850), .B(pin_io[53]), .O(pin_io_out_53));
    BB pin_io_pad_54 (.I(GND_net), .T(VCC_net), .B(pin_io[54]), .O(pin_io_out_54));   // c:/s_links/sources/slot_cards/shutter_4.v(70[8:14])
    BB pin_io_pad_55 (.I(n26523), .T(n26579), .B(pin_io[55]), .O(pin_io_out_55));
    BB pin_io_pad_56 (.I(n2_adj_7965), .T(n8661), .B(pin_io[56]), .O(pin_io_out_56));
    BB pin_io_pad_58 (.I(GND_net), .T(VCC_net), .B(pin_io[58]), .O(pin_io_out_58));   // c:/s_links/sources/slot_cards/shutter_4.v(73[8:14])
    BB pin_io_pad_59 (.I(n1_adj_8157), .T(n8840), .B(pin_io[59]), .O(pin_io_out_59));
    BB pin_io_pad_62 (.I(GND_net), .T(VCC_net), .B(pin_io[62]), .O(pin_io_out_62));   // c:/s_links/sources/slot_cards/shutter_4.v(68[8:14])
    BB pin_io_pad_63 (.I(n2_adj_8155), .T(n8836), .B(pin_io[63]), .O(pin_io_out_63));
    BB pin_io_pad_64 (.I(GND_net), .T(VCC_net), .B(pin_io[64]), .O(pin_io_out_64));   // c:/s_links/sources/slot_cards/shutter_4.v(70[8:14])
    BB pin_io_pad_65 (.I(n26521), .T(n28813), .B(pin_io[65]), .O(pin_io_out_65));
    BB pin_io_pad_66 (.I(n2_adj_7620), .T(n8633), .B(pin_io[66]), .O(pin_io_out_66));
    BB pin_io_pad_68 (.I(GND_net), .T(VCC_net), .B(pin_io[68]), .O(pin_io_out_68));   // c:/s_links/sources/slot_cards/shutter_4.v(73[8:14])
    LUT4 i22851_2_lut (.A(n19351), .B(resetn_c), .Z(clk_1MHz_enable_91)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i22851_2_lut.init = 16'h7777;
    LUT4 i22697_2_lut (.A(n19391), .B(resetn_c), .Z(clk_1MHz_enable_40)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i22697_2_lut.init = 16'h7777;
    \io(DEV_ID=3,UART_ADDRESS_WIDTH=4)  \io_ins_3..u_io  (.mode(mode_adj_8131), 
            .clk(clk), .clk_enable_201(clk_enable_201), .n29239(n29239), 
            .\spi_data_r[0] (spi_data_r[0])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(464[3] 496[2])
    \shutter(DEV_ID=3,UART_ADDRESS_WIDTH=4)  \shutter_ins_3..u_shutter  (.\mode[1] (n29783[1]), 
            .\mode[2] (n29783[2]), .n29225(n29225), .\quad_homing[1] (quad_homing_adj_8343[1]), 
            .n27632(n27632), .n26969(n26969), .n13052(n13052), .pin_io_out_34(pin_io_out_34), 
            .\pin_intrpt[11] (pin_intrpt[11]), .pin_io_out_32(pin_io_out_32), 
            .\pin_intrpt[9] (pin_intrpt[9]), .reset_r(reset_r_adj_7981), 
            .n1(n1_adj_8167), .\cs_decoded[6] (cs_decoded[6]), .n2(n2_adj_7957), 
            .pin_io_out_33(pin_io_out_33), .\pin_intrpt[10] (pin_intrpt[10]), 
            .mode(mode_adj_8139), .clk(clk), .clk_enable_171(clk_enable_171), 
            .n29239(n29239), .\spi_data_r[0] (spi_data_r[0])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(508[3] 540[2])
    \shutter(DEV_ID=2,UART_ADDRESS_WIDTH=4)  \shutter_ins_2..u_shutter  (.\mode[1] (n29782[1]), 
            .\mode[2] (n29782[2]), .n29233(n29233), .pin_io_out_22(pin_io_out_22), 
            .\pin_intrpt[6] (pin_intrpt[6]), .reset_r(reset_r_adj_7975), 
            .n1(n1_adj_8171), .\cs_decoded[4] (cs_decoded[4]), .n2(n2_adj_7964), 
            .pin_io_out_24(pin_io_out_24), .\mode[2]_derived_32 (mode_2_derived_32_adj_8013), 
            .pin_io_out_23(pin_io_out_23), .\pin_intrpt[7] (pin_intrpt[7]), 
            .mode(mode_adj_8138), .clk(clk), .clk_enable_176(clk_enable_176), 
            .n29239(n29239), .\spi_data_r[0] (spi_data_r[0]), .n29194(n29194), 
            .n29193(n29193), .n29303(n29303), .n27480(n27480)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(508[3] 540[2])
    \shutter(DEV_ID=4,UART_ADDRESS_WIDTH=4)  \shutter_ins_4..u_shutter  (.\mode[1] (n29784[1]), 
            .\mode[2] (n29784[2]), .n29224(n29224), .pin_io_out_44(pin_io_out_44), 
            .\pin_intrpt[14] (pin_intrpt[14]), .pin_io_out_42(pin_io_out_42), 
            .\pin_intrpt[12] (pin_intrpt[12]), .reset_r(reset_r_adj_8017), 
            .n1(n1_adj_8164), .\cs_decoded[8] (cs_decoded[8]), .n2(n2), 
            .pin_io_out_43(pin_io_out_43), .\pin_intrpt[13] (pin_intrpt[13]), 
            .mode(mode_adj_8140), .clk(clk), .clk_enable_169(clk_enable_169), 
            .n29239(n29239), .\spi_data_r[0] (spi_data_r[0])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(508[3] 540[2])
    \io(DEV_ID=4,UART_ADDRESS_WIDTH=4)  \io_ins_4..u_io  (.mode(mode_adj_8132), 
            .clk(clk), .clk_enable_166(clk_enable_166), .n29239(n29239), 
            .\spi_data_r[0] (spi_data_r[0])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(464[3] 496[2])
    \quad_decoder(DEV_ID=6)  \quad_ins_6..u_quad_decoder  (.quad_count({quad_count_adj_8521}), 
            .clk_1MHz(clk_1MHz), .\spi_data_out_r_39__N_2338[0] (spi_data_out_r_39__N_2338[0]), 
            .clk(clk), .\spi_data_out_r_39__N_2483[0] (spi_data_out_r_39__N_2483[0]), 
            .\quad_b[6] (quad_b[6]), .quad_buffer({quad_buffer_adj_8522}), 
            .\pin_intrpt[20] (pin_intrpt[20]), .n29239(n29239), .clk_enable_76(clk_enable_76), 
            .\spi_data_r[31] (spi_data_r[31]), .\spi_data_r[30] (spi_data_r[30]), 
            .\spi_data_r[29] (spi_data_r[29]), .\spi_data_r[28] (spi_data_r[28]), 
            .\spi_data_r[27] (spi_data_r[27]), .\spi_data_r[26] (spi_data_r[26]), 
            .\spi_data_r[25] (spi_data_r[25]), .\spi_data_r[24] (spi_data_r[24]), 
            .\spi_data_r[23] (spi_data_r[23]), .\spi_data_r[22] (spi_data_r[22]), 
            .\spi_data_r[21] (spi_data_r[21]), .\spi_data_r[20] (spi_data_r[20]), 
            .\spi_data_r[19] (spi_data_r[19]), .\spi_data_r[0] (spi_data_r[0]), 
            .\spi_data_r[18] (spi_data_r[18]), .\spi_data_r[17] (spi_data_r[17]), 
            .\spi_data_r[16] (spi_data_r[16]), .\spi_data_r[15] (spi_data_r[15]), 
            .\spi_data_r[14] (spi_data_r[14]), .\spi_data_r[13] (spi_data_r[13]), 
            .\spi_data_r[12] (spi_data_r[12]), .\spi_data_r[11] (spi_data_r[11]), 
            .\spi_data_r[10] (spi_data_r[10]), .\spi_data_r[9] (spi_data_r[9]), 
            .\spi_data_r[8] (spi_data_r[8]), .\spi_data_r[7] (spi_data_r[7]), 
            .\spi_data_r[6] (spi_data_r[6]), .\spi_data_r[5] (spi_data_r[5]), 
            .\spi_data_r[4] (spi_data_r[4]), .\spi_data_r[3] (spi_data_r[3]), 
            .\spi_data_r[2] (spi_data_r[2]), .\spi_data_r[1] (spi_data_r[1]), 
            .clk_enable_499(clk_enable_499), .n29762(n29762), .resetn_c(resetn_c), 
            .GND_net(GND_net), .spi_data_out_r_39__N_2378(spi_data_out_r_39__N_2378), 
            .spi_data_out_r_39__N_2566(spi_data_out_r_39__N_2566), .quad_set_complete(quad_set_complete_adj_7891), 
            .\quad_a[6] (quad_a[6]), .\spi_data_out_r_39__N_2338[31] (spi_data_out_r_39__N_2338[31]), 
            .\spi_data_out_r_39__N_2483[31] (spi_data_out_r_39__N_2483[31]), 
            .\spi_data_out_r_39__N_2338[30] (spi_data_out_r_39__N_2338[30]), 
            .\spi_data_out_r_39__N_2483[30] (spi_data_out_r_39__N_2483[30]), 
            .\spi_data_out_r_39__N_2338[29] (spi_data_out_r_39__N_2338[29]), 
            .\spi_data_out_r_39__N_2483[29] (spi_data_out_r_39__N_2483[29]), 
            .\spi_data_out_r_39__N_2338[28] (spi_data_out_r_39__N_2338[28]), 
            .\spi_data_out_r_39__N_2483[28] (spi_data_out_r_39__N_2483[28]), 
            .\spi_data_out_r_39__N_2338[27] (spi_data_out_r_39__N_2338[27]), 
            .\spi_data_out_r_39__N_2483[27] (spi_data_out_r_39__N_2483[27]), 
            .\spi_data_out_r_39__N_2338[26] (spi_data_out_r_39__N_2338[26]), 
            .\spi_data_out_r_39__N_2483[26] (spi_data_out_r_39__N_2483[26]), 
            .\spi_data_out_r_39__N_2338[25] (spi_data_out_r_39__N_2338[25]), 
            .\spi_data_out_r_39__N_2483[25] (spi_data_out_r_39__N_2483[25]), 
            .\spi_data_out_r_39__N_2338[24] (spi_data_out_r_39__N_2338[24]), 
            .\spi_data_out_r_39__N_2483[24] (spi_data_out_r_39__N_2483[24]), 
            .\spi_data_out_r_39__N_2338[23] (spi_data_out_r_39__N_2338[23]), 
            .\spi_data_out_r_39__N_2483[23] (spi_data_out_r_39__N_2483[23]), 
            .\spi_data_out_r_39__N_2338[22] (spi_data_out_r_39__N_2338[22]), 
            .\spi_data_out_r_39__N_2483[22] (spi_data_out_r_39__N_2483[22]), 
            .\spi_data_out_r_39__N_2338[21] (spi_data_out_r_39__N_2338[21]), 
            .\spi_data_out_r_39__N_2483[21] (spi_data_out_r_39__N_2483[21]), 
            .\spi_data_out_r_39__N_2338[20] (spi_data_out_r_39__N_2338[20]), 
            .\spi_data_out_r_39__N_2483[20] (spi_data_out_r_39__N_2483[20]), 
            .\spi_data_out_r_39__N_2338[19] (spi_data_out_r_39__N_2338[19]), 
            .\spi_data_out_r_39__N_2483[19] (spi_data_out_r_39__N_2483[19]), 
            .\spi_data_out_r_39__N_2338[18] (spi_data_out_r_39__N_2338[18]), 
            .\spi_data_out_r_39__N_2483[18] (spi_data_out_r_39__N_2483[18]), 
            .\spi_data_out_r_39__N_2338[17] (spi_data_out_r_39__N_2338[17]), 
            .\spi_data_out_r_39__N_2483[17] (spi_data_out_r_39__N_2483[17]), 
            .\spi_data_out_r_39__N_2338[16] (spi_data_out_r_39__N_2338[16]), 
            .\spi_data_out_r_39__N_2483[16] (spi_data_out_r_39__N_2483[16]), 
            .\spi_data_out_r_39__N_2338[15] (spi_data_out_r_39__N_2338[15]), 
            .\spi_data_out_r_39__N_2483[15] (spi_data_out_r_39__N_2483[15]), 
            .\spi_data_out_r_39__N_2338[14] (spi_data_out_r_39__N_2338[14]), 
            .\spi_data_out_r_39__N_2483[14] (spi_data_out_r_39__N_2483[14]), 
            .\spi_data_out_r_39__N_2338[13] (spi_data_out_r_39__N_2338[13]), 
            .\spi_data_out_r_39__N_2483[13] (spi_data_out_r_39__N_2483[13]), 
            .\spi_data_out_r_39__N_2338[12] (spi_data_out_r_39__N_2338[12]), 
            .\spi_data_out_r_39__N_2483[12] (spi_data_out_r_39__N_2483[12]), 
            .\spi_data_out_r_39__N_2338[11] (spi_data_out_r_39__N_2338[11]), 
            .\spi_data_out_r_39__N_2483[11] (spi_data_out_r_39__N_2483[11]), 
            .\spi_data_out_r_39__N_2338[10] (spi_data_out_r_39__N_2338[10]), 
            .\spi_data_out_r_39__N_2483[10] (spi_data_out_r_39__N_2483[10]), 
            .\spi_data_out_r_39__N_2338[9] (spi_data_out_r_39__N_2338[9]), 
            .\spi_data_out_r_39__N_2483[9] (spi_data_out_r_39__N_2483[9]), 
            .\spi_data_out_r_39__N_2338[8] (spi_data_out_r_39__N_2338[8]), 
            .\spi_data_out_r_39__N_2483[8] (spi_data_out_r_39__N_2483[8]), 
            .\spi_data_out_r_39__N_2338[7] (spi_data_out_r_39__N_2338[7]), 
            .\spi_data_out_r_39__N_2483[7] (spi_data_out_r_39__N_2483[7]), 
            .\spi_data_out_r_39__N_2338[6] (spi_data_out_r_39__N_2338[6]), 
            .\spi_data_out_r_39__N_2483[6] (spi_data_out_r_39__N_2483[6]), 
            .\spi_data_out_r_39__N_2338[5] (spi_data_out_r_39__N_2338[5]), 
            .\spi_data_out_r_39__N_2483[5] (spi_data_out_r_39__N_2483[5]), 
            .\spi_data_out_r_39__N_2338[4] (spi_data_out_r_39__N_2338[4]), 
            .\spi_data_out_r_39__N_2483[4] (spi_data_out_r_39__N_2483[4]), 
            .\spi_data_out_r_39__N_2338[3] (spi_data_out_r_39__N_2338[3]), 
            .\spi_data_out_r_39__N_2483[3] (spi_data_out_r_39__N_2483[3]), 
            .\spi_data_out_r_39__N_2338[2] (spi_data_out_r_39__N_2338[2]), 
            .\spi_data_out_r_39__N_2483[2] (spi_data_out_r_39__N_2483[2]), 
            .\spi_data_out_r_39__N_2338[1] (spi_data_out_r_39__N_2338[1]), 
            .\spi_data_out_r_39__N_2483[1] (spi_data_out_r_39__N_2483[1]), 
            .pin_io_out_64(pin_io_out_64), .n29267(n29267), .clk_enable_520(clk_enable_520), 
            .n29092(n29092)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(272[3] 293[2])
    \io(DEV_ID=5,UART_ADDRESS_WIDTH=4)  \io_ins_5..u_io  (.mode(mode_adj_8133), 
            .clk(clk), .clk_enable_182(clk_enable_182), .n29239(n29239), 
            .\spi_data_r[0] (spi_data_r[0])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(464[3] 496[2])
    \io(UART_ADDRESS_WIDTH=4)  \io_ins_0..u_io  (.mode(mode_adj_8128), .clk(clk), 
            .clk_enable_167(clk_enable_167), .n29239(n29239), .\spi_data_r[0] (spi_data_r[0]), 
            .\spi_cmd_r[2] (spi_cmd_r[2]), .\spi_addr_r[2] (spi_addr_r[2]), 
            .n29256(n29256), .n29101(n29101), .resetn_c(resetn_c), .clk_enable_178(clk_enable_178), 
            .n19233(n19233), .\spi_addr_r[0] (spi_addr_r[0]), .\spi_cmd_r[1] (spi_cmd_r[1]), 
            .n29288(n29288), .n65(n65_adj_8152), .n29110(n29110), .\spi_cmd_r[0] (spi_cmd_r[0]), 
            .n27058(n27058), .n13074(n13074), .n29213(n29213), .\spi_cmd[1] (spi_cmd[1]), 
            .\spi_addr_r[3] (spi_addr_r[3]), .spi_sdo_valid_N_297(spi_sdo_valid_N_297), 
            .spi_sdo_valid_N_296(spi_sdo_valid_N_296), .\spi_cmd[2] (spi_cmd[2]), 
            .\spi_cmd[15] (spi_cmd[15]), .n29761(n29761), .n19084(n19084), 
            .n27618(n27618), .n31(n31_adj_8153), .\spi_cmd[4] (spi_cmd[4]), 
            .n29144(n29144), .n29182(n29182), .n29169(n29169), .n29114(n29114), 
            .\spi_addr_r[1] (spi_addr_r[1]), .n29214(n29214), .n29105(n29105), 
            .n29211(n29211), .n27225(n27225), .n29120(n29120)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(464[3] 496[2])
    \io(DEV_ID=2,UART_ADDRESS_WIDTH=4)  \io_ins_2..u_io  (.mode(mode_adj_8130), 
            .clk(clk), .clk_enable_202(clk_enable_202), .n29239(n29239), 
            .\spi_data_r[0] (spi_data_r[0])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(464[3] 496[2])
    \io(DEV_ID=1,UART_ADDRESS_WIDTH=4)  \io_ins_1..u_io  (.mode(mode_adj_8129), 
            .clk(clk), .clk_enable_197(clk_enable_197), .n29239(n29239), 
            .\spi_data_r[0] (spi_data_r[0])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(464[3] 496[2])
    LUT4 i22777_2_lut (.A(n19381), .B(resetn_c), .Z(clk_1MHz_enable_66)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i22777_2_lut.init = 16'h7777;
    \servo(DEV_ID=3,UART_ADDRESS_WIDTH=4)  \servo_ins_3..u_servo  (.mode(mode_adj_8124), 
            .clk(clk), .clk_enable_180(clk_enable_180), .n29239(n29239), 
            .n29762(n29762), .n29196(n29196), .C_5_c_c(C_5_c_c), .n29225(n29225), 
            .n8720(n8720)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(418[3] 453[2])
    \servo(DEV_ID=1,UART_ADDRESS_WIDTH=4)  \servo_ins_1..u_servo  (.mode(mode_adj_8122), 
            .clk(clk), .clk_enable_184(clk_enable_184), .n29239(n29239), 
            .n29762(n29762), .n29202(n29202), .C_5_c_c(C_5_c_c), .n29237(n29237), 
            .n8777(n8777)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(418[3] 453[2])
    \servo(DEV_ID=2,UART_ADDRESS_WIDTH=4)  \servo_ins_2..u_servo  (.mode(mode_adj_8123), 
            .clk(clk), .clk_enable_181(clk_enable_181), .n29239(n29239), 
            .n29762(n29762), .n29194(n29194), .C_5_c_c(C_5_c_c), .n29233(n29233), 
            .n8749(n8749)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(418[3] 453[2])
    \servo(DEV_ID=5,UART_ADDRESS_WIDTH=4)  \servo_ins_5..u_servo  (.mode(mode_adj_8126), 
            .clk(clk), .clk_enable_175(clk_enable_175), .n29239(n29239), 
            .n29762(n29762), .n29199(n29199), .C_5_c_c(C_5_c_c), .n29220(n29220), 
            .n8661(n8661)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(418[3] 453[2])
    \servo(UART_ADDRESS_WIDTH=4)  \servo_ins_0..u_servo  (.mode(mode), .n29160(n29160), 
            .C_5_c_c(C_5_c_c), .n29260(n29260), .n8805(n8805), .clk(clk), 
            .clk_enable_186(clk_enable_186), .n29239(n29239), .n29762(n29762)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(418[3] 453[2])
    \servo(DEV_ID=4,UART_ADDRESS_WIDTH=4)  \servo_ins_4..u_servo  (.mode(mode_adj_8125), 
            .clk(clk), .clk_enable_178(clk_enable_178), .n29239(n29239), 
            .n29762(n29762), .n29204(n29204), .C_5_c_c(C_5_c_c), .n29224(n29224), 
            .n8689(n8689)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(418[3] 453[2])
    \otm_dac(DEV_ID=3)  u_otm_dac (.NSL(NSL), .n29317(n29317), .mode(mode_adj_8143), 
            .n8717(n8717), .clk(clk), .clk_enable_193(clk_enable_193), 
            .n29239(n29239), .\spi_data_r[0] (spi_data_r[0]), .clk_enable_204(clk_enable_204), 
            .n29214(n29214), .n29127(n29127), .n27259(n27259), .\spi_addr_r[1] (spi_addr_r[1]), 
            .n29084(n29084), .n29254(n29254), .n27286(n27286), .reset_r_N_4813(reset_r_N_4813), 
            .n29162(n29162), .n29085(n29085)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(577[3] 595[2])
    LUT4 i22601_2_lut (.A(n19337), .B(resetn_c), .Z(clk_1MHz_enable_55)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i22601_2_lut.init = 16'h7777;
    \shutter(DEV_ID=1,UART_ADDRESS_WIDTH=4)  \shutter_ins_1..u_shutter  (.mode_adj_554({n29781}), 
            .n29237(n29237), .\quad_homing[1] (quad_homing_adj_8225[1]), 
            .n27636(n27636), .n26963(n26963), .n12716(n12716), .pin_io_out_14(pin_io_out_14), 
            .\pin_intrpt[5] (pin_intrpt[5]), .pin_io_out_12(pin_io_out_12), 
            .\pin_intrpt[3] (pin_intrpt[3]), .reset_r(reset_r_adj_7969), 
            .n1(n1_adj_8175), .\cs_decoded[2] (cs_decoded[2]), .n2(n2_adj_7971), 
            .n29198(n29198), .pin_io_out_13(pin_io_out_13), .\pin_intrpt[4] (pin_intrpt[4]), 
            .mode(mode_adj_8137), .clk(clk), .clk_enable_179(clk_enable_179), 
            .n29239(n29239), .\spi_data_r[0] (spi_data_r[0]), .n8898(n8898)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(508[3] 540[2])
    \peizo_elliptec(DEV_ID=7,UART_ADDRESS_WIDTH=4)  u_peizo_elliptec (.clk(clk), 
            .clk_enable_194(clk_enable_194), .n29239(n29239), .\spi_data_r[0] (spi_data_r[0]), 
            .C_1_c_0(C_1_c_0), .n29313(n29313), .C_2_c_1(C_2_c_1), .tx_N_6443(tx_N_6443)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(602[3] 622[2])
    LUT4 i2732_4_lut (.A(spi_cmd_valid), .B(n29247), .C(spi_addr_valid), 
         .D(spi_data_valid), .Z(clk_enable_524)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;
    defparam i2732_4_lut.init = 16'hcdcc;
    BB pin_io_pad_69 (.I(n1), .T(n8826), .B(pin_io[69]), .O(pin_io_out_69));
    \shutter(UART_ADDRESS_WIDTH=4)  \shutter_ins_0..u_shutter  (.mode(mode_adj_8135), 
            .clk(clk), .clk_enable_189(clk_enable_189), .n29239(n29239), 
            .\spi_data_r[0] (spi_data_r[0]), .\mode[1] (n29780[1]), .\mode[2] (n29780[2]), 
            .n29260(n29260), .\quad_homing[0] (quad_homing[0]), .pin_io_out_4(pin_io_out_4), 
            .n5(n5_adj_8136), .pin_io_out_2(pin_io_out_2), .\pin_intrpt[0] (pin_intrpt[0]), 
            .reset_r(reset_r), .n1(n1_adj_8179), .\cs_decoded[0] (cs_decoded[0]), 
            .n2(n2_adj_7977), .\mode[2]_derived_32 (mode_2_derived_32), 
            .pin_io_out_3(pin_io_out_3), .\pin_intrpt[1] (pin_intrpt[1]), 
            .n29160(n29160), .mode_adj_553(mode_adj_8128), .n29201(n29201), 
            .n31(n31_adj_8085), .n27471(n27471), .n29089(n29089), .n29254(n29254), 
            .n29083(n29083), .resetn_c(resetn_c), .clk_enable_198(clk_enable_198), 
            .n29214(n29214), .n29118(n29118), .\spi_addr_r[1] (spi_addr_r[1]), 
            .n27256(n27256), .reset_r_N_4474(reset_r_N_4474), .n19084(n19084), 
            .\spi_cmd_r[1] (spi_cmd_r[1]), .\spi_cmd_r[3] (spi_cmd_r[3]), 
            .n29082(n29082), .n29182(n29182), .\spi_cmd_r[0] (spi_cmd_r[0]), 
            .n29130(n29130), .n65(n65_adj_8152), .n27(n27), .\spi_addr_r[2] (spi_addr_r[2]), 
            .n27283(n27283), .clk_enable_164(clk_enable_164), .n29174(n29174), 
            .n29127(n29127), .n27285(n27285), .n29104(n29104), .n29251(n29251), 
            .n29256(n29256), .n29102(n29102), .n19233(n19233), .n29100(n29100), 
            .n29096(n29096), .n13074(n13074), .clk_enable_173(clk_enable_173)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(508[3] 540[2])
    LUT4 i22823_2_lut (.A(n19371), .B(resetn_c), .Z(clk_1MHz_enable_182)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i22823_2_lut.init = 16'h7777;
    \piezo(DEV_ID=1,UART_ADDRESS_WIDTH=4)  \piezo_ins_1..u_piezo  (.mode(mode_adj_8145), 
            .clk(clk), .clk_enable_187(clk_enable_187), .n29239(n29239), 
            .\spi_data_r[0] (spi_data_r[0]), .n29282(n29282), .n29284(n29284), 
            .n29237(n29237), .mode_adj_552({n29781}), .OW_ID_N_4464(OW_ID_N_4464), 
            .C_1_c_0(C_1_c_0), .C_2_c_1(C_2_c_1), .mode_adj_549(mode_adj_8126), 
            .n29313(n29313), .n29158(n29158), .mode_adj_550(mode_adj_8122), 
            .n29157(n29157), .n13(n13_adj_8151), .n27483(n27483), .\cs_decoded[3] (cs_decoded[3]), 
            .n2(n2_adj_8174), .n8908(n8908), .digital_output_r(digital_output_r_adj_7970), 
            .n26533(n26533), .OW_ID_N_4462(OW_ID_N_4462), .C_5_c_c(C_5_c_c), 
            .n29202(n29202), .n13615(n13615), .mode_adj_551(mode_adj_8129), 
            .n29306(n29306), .n29315(n29315), .n8795(n8795)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(632[3] 661[2])
    \piezo(UART_ADDRESS_WIDTH=4)  \piezo_ins_0..u_piezo  (.mode(mode_adj_8144), 
            .clk(clk), .clk_enable_192(clk_enable_192), .n29239(n29239), 
            .\spi_data_r[0] (spi_data_r[0]), .\spi_cmd_r[3] (spi_cmd_r[3]), 
            .n29251(n29251), .\spi_addr_r[1] (spi_addr_r[1]), .n29214(n29214), 
            .n29124(n29124), .mode_adj_548({n29780}), .digital_output_r(digital_output_r), 
            .n26535(n26535), .n26561(n26561), .n27(n27), .\spi_addr_r[2] (spi_addr_r[2]), 
            .n29161(n29161), .n29169(n29169), .n29216(n29216), .n27225(n27225), 
            .\spi_addr_r[0] (spi_addr_r[0]), .n19084(n19084), .n29286(n29286), 
            .n29123(n29123), .n29287(n29287), .n29101(n29101), .\cs_decoded[1] (cs_decoded[1]), 
            .n2(n2_adj_8178), .n8922(n8922), .C_5_c_c(C_5_c_c), .n22(n22), 
            .C_4_c_3(C_4_c_3), .n29200(n29200), .n3(n3_adj_7963), .n29307(n29307), 
            .\spi_cmd_r[1] (spi_cmd_r[1]), .n27240(n27240), .mode_adj_547(mode_adj_8128), 
            .n29309(n29309), .\spi_cmd_r[2] (spi_cmd_r[2]), .n29288(n29288), 
            .n65(n65), .n27234(n27234)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(632[3] 661[2])
    LUT4 i22684_2_lut (.A(n19401), .B(resetn_c), .Z(clk_1MHz_enable_367)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i22684_2_lut.init = 16'h7777;
    \piezo(DEV_ID=2,UART_ADDRESS_WIDTH=4)  \piezo_ins_2..u_piezo  (.mode(mode_adj_8146), 
            .clk(clk), .clk_enable_185(clk_enable_185), .n29239(n29239), 
            .n29762(n29762), .\cs_decoded[5] (cs_decoded[5]), .n2(n2_adj_8170), 
            .n8894(n8894), .mode_adj_546({n29782}), .digital_output_r(digital_output_r_adj_7976), 
            .n26531(n26531), .n26549(n26549), .n27590(n27590), .C_2_c_1(C_2_c_1), 
            .C_1_c_0(C_1_c_0), .n22(n22_adj_7754), .n8884(n8884)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(632[3] 661[2])
    \piezo(DEV_ID=3,UART_ADDRESS_WIDTH=4)  \piezo_ins_3..u_piezo  (.mode(mode_adj_8147), 
            .clk(clk), .clk_enable_183(clk_enable_183), .n29239(n29239), 
            .n29762(n29762), .n29203(n29203), .n29300(n29300), .mode_adj_544(mode_adj_8139), 
            .pin_io_out_35(pin_io_out_35), .n26972(n26972), .\cs_decoded[7] (cs_decoded[7]), 
            .n2(n2_adj_8166), .n8880(n8880), .mode_adj_545({n29783}), 
            .digital_output_r(digital_output_r_adj_7982), .n26529(n26529), 
            .n26565(n26565), .n27590(n27590), .C_1_c_0(C_1_c_0), .C_2_c_1(C_2_c_1), 
            .n29149(n29149), .n8870(n8870)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(632[3] 661[2])
    \piezo(DEV_ID=4,UART_ADDRESS_WIDTH=4)  \piezo_ins_4..u_piezo  (.mode(mode_adj_8148), 
            .clk(clk), .clk_enable_177(clk_enable_177), .n29239(n29239), 
            .n29762(n29762), .mode_adj_543({n29784}), .digital_output_r(digital_output_r_adj_8018), 
            .n26525(n26525), .C_4_c_3(C_4_c_3), .n29200(n29200), .pin_io_out_6(pin_io_out_6), 
            .mode_adj_539(mode), .n7(n7), .C_3_c_2(C_3_c_2), .n29132(n29132), 
            .C_1_c_0(C_1_c_0), .C_2_c_1(C_2_c_1), .n29160(n29160), .mode_adj_540(mode_adj_8125), 
            .n29284(n29284), .n29150(n29150), .n29196(n29196), .n29202(n29202), 
            .n29204(n29204), .C_5_c_c(C_5_c_c), .n27590(n27590), .n29194(n29194), 
            .OW_ID_N_5482(OW_ID_N_5482), .mode_adj_541(mode_adj_8132), .n27189(n27189), 
            .mode_adj_542(mode_adj_8140), .\cs_decoded[9] (cs_decoded[9]), 
            .n2(n2_adj_8163), .n8864(n8864), .n26569(n26569), .n8854(n8854)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(632[3] 661[2])
    \intrpt_ctrl(DEV_ID=5)  \intrpt_ins_5..u_intrpt_ctrl  (.\spi_data_out_r_39__N_2927[0] (spi_data_out_r_39__N_2927[0]), 
            .clk(clk), .\pin_intrpt[15] (pin_intrpt[15]), .n29239(n29239), 
            .clear_intrpt(clear_intrpt_adj_7961), .clear_intrpt_N_2994(clear_intrpt_N_2994), 
            .intrpt_out_c_5(intrpt_out_c_5), .intrpt_out_N_2990(intrpt_out_N_2990), 
            .n29757(n29757), .\spi_data_out_r_39__N_2927[2] (spi_data_out_r_39__N_2927[2]), 
            .\mode[2]_derived_32 (mode_2_derived_32_adj_8049), .\spi_data_out_r_39__N_2927[1] (spi_data_out_r_39__N_2927[1]), 
            .\pin_intrpt[16] (pin_intrpt[16])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(304[3] 325[2])
    \shutter(DEV_ID=6,UART_ADDRESS_WIDTH=4)  \shutter_ins_6..u_shutter  (.mode(mode_adj_8142), 
            .clk(clk), .clk_enable_32(clk_enable_32), .n29239(n29239), 
            .\spi_data_r[0] (spi_data_r[0]), .mode_adj_538({n29786}), .n29267(n29267), 
            .pin_io_out_64(pin_io_out_64), .\pin_intrpt[20] (pin_intrpt[20]), 
            .pin_io_out_62(pin_io_out_62), .\pin_intrpt[18] (pin_intrpt[18]), 
            .pin_io_out_63(pin_io_out_63), .\pin_intrpt[19] (pin_intrpt[19]), 
            .reset_r(reset_r_adj_8089), .n1(n1_adj_8156), .\cs_decoded[12] (cs_decoded[12]), 
            .n2(n2_adj_7620), .n29190(n29190), .n8826(n8826)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(508[3] 540[2])
    \shutter(DEV_ID=5,UART_ADDRESS_WIDTH=4)  \shutter_ins_5..u_shutter  (.\mode[1] (n29785[1]), 
            .\mode[2] (n29785[2]), .n29220(n29220), .\quad_homing[0] (quad_homing_adj_8461[0]), 
            .pin_io_out_54(pin_io_out_54), .n27657(n27657), .pin_io_out_52(pin_io_out_52), 
            .\pin_intrpt[15] (pin_intrpt[15]), .reset_r(reset_r_adj_8053), 
            .n1(n1_adj_8160), .\cs_decoded[10] (cs_decoded[10]), .n2(n2_adj_7965), 
            .\mode[2]_derived_32 (mode_2_derived_32_adj_8049), .pin_io_out_53(pin_io_out_53), 
            .\pin_intrpt[16] (pin_intrpt[16]), .mode(mode_adj_8141), .clk(clk), 
            .clk_enable_172(clk_enable_172), .n29239(n29239), .\spi_data_r[0] (spi_data_r[0])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(508[3] 540[2])
    \io(DEV_ID=6,UART_ADDRESS_WIDTH=4)  \io_ins_6..u_io  (.mode(mode_adj_8134), 
            .clk(clk), .clk_enable_191(clk_enable_191), .n29239(n29239), 
            .\spi_data_r[0] (spi_data_r[0])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(464[3] 496[2])
    \status_led(DEV_ID=9)  u_status_led (.clk(clk), .resetn_c(resetn_c), 
            .clk_enable_303(clk_enable_303), .n29239(n29239), .\spi_data_r[0] (spi_data_r[0]), 
            .GND_net(GND_net), .\spi_data_out_r_39__N_770[0] (spi_data_out_r_39__N_770[0]), 
            .spi_data_out_r_39__N_810(spi_data_out_r_39__N_810), .EM_STOP(EM_STOP), 
            .led_sw_c(led_sw_c), .\spi_cmd_r[8] (spi_cmd_r[8]), .n13265(n13265), 
            .\spi_cmd_r[14] (spi_cmd_r[14]), .\spi_cmd_r[11] (spi_cmd_r[11]), 
            .\spi_cmd_r[9] (spi_cmd_r[9]), .\spi_cmd_r[13] (spi_cmd_r[13]), 
            .\spi_cmd_r[7] (spi_cmd_r[7]), .\spi_cmd_r[10] (spi_cmd_r[10]), 
            .spi_data_valid_r(spi_data_valid_r), .\spi_cmd_r[12] (spi_cmd_r[12]), 
            .\spi_cmd_r[6] (spi_cmd_r[6]), .\spi_cmd_r[15] (spi_cmd_r[15]), 
            .\spi_data_r[11] (spi_data_r[11]), .\spi_data_r[10] (spi_data_r[10]), 
            .\spi_data_r[9] (spi_data_r[9]), .\spi_data_r[8] (spi_data_r[8]), 
            .\spi_data_r[7] (spi_data_r[7]), .\spi_data_r[6] (spi_data_r[6]), 
            .\spi_data_r[5] (spi_data_r[5]), .\spi_data_r[4] (spi_data_r[4]), 
            .\spi_data_r[3] (spi_data_r[3]), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[1] (spi_data_r[1]), .n6(n6), .\spi_addr[3] (spi_addr[3]), 
            .n27465(n27465), .\spi_cmd[1] (spi_cmd[1]), .\spi_addr[0] (spi_addr[0]), 
            .n13489(n13489), .n26928(n26928)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(228[3] 245[2])
    \intrpt_ctrl(DEV_ID=4)  \intrpt_ins_4..u_intrpt_ctrl  (.\spi_data_out_r_39__N_2856[0] (spi_data_out_r_39__N_2856[0]), 
            .clk(clk), .\pin_intrpt[12] (pin_intrpt[12]), .n29239(n29239), 
            .clear_intrpt(clear_intrpt_adj_7960), .clear_intrpt_N_2923(clear_intrpt_N_2923), 
            .intrpt_out_c_4(intrpt_out_c_4), .intrpt_out_N_2919(intrpt_out_N_2919), 
            .n29757(n29757), .\spi_data_out_r_39__N_2856[2] (spi_data_out_r_39__N_2856[2]), 
            .\pin_intrpt[14] (pin_intrpt[14]), .\spi_data_out_r_39__N_2856[1] (spi_data_out_r_39__N_2856[1]), 
            .\pin_intrpt[13] (pin_intrpt[13])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(304[3] 325[2])
    \intrpt_ctrl(DEV_ID=3)  \intrpt_ins_3..u_intrpt_ctrl  (.clk(clk), .n29239(n29239), 
            .\spi_data_out_r_39__N_2785[0] (spi_data_out_r_39__N_2785[0]), 
            .\pin_intrpt[9] (pin_intrpt[9]), .clear_intrpt(clear_intrpt_adj_7959), 
            .clear_intrpt_N_2852(clear_intrpt_N_2852), .intrpt_out_c_3(intrpt_out_c_3), 
            .intrpt_out_N_2848(intrpt_out_N_2848), .n29757(n29757), .\spi_data_out_r_39__N_2785[2] (spi_data_out_r_39__N_2785[2]), 
            .\pin_intrpt[11] (pin_intrpt[11]), .\spi_data_out_r_39__N_2785[1] (spi_data_out_r_39__N_2785[1]), 
            .\pin_intrpt[10] (pin_intrpt[10])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(304[3] 325[2])
    \intrpt_ctrl(DEV_ID=2)  \intrpt_ins_2..u_intrpt_ctrl  (.clk(clk), .n29239(n29239), 
            .\spi_data_out_r_39__N_2714[0] (spi_data_out_r_39__N_2714[0]), 
            .\pin_intrpt[6] (pin_intrpt[6]), .intrpt_out_c_2(intrpt_out_c_2), 
            .intrpt_out_N_2777(intrpt_out_N_2777), .n29757(n29757), .clear_intrpt(clear_intrpt_adj_7958), 
            .clear_intrpt_N_2781(clear_intrpt_N_2781), .\spi_data_out_r_39__N_2714[2] (spi_data_out_r_39__N_2714[2]), 
            .\mode[2]_derived_32 (mode_2_derived_32_adj_8013), .\spi_data_out_r_39__N_2714[1] (spi_data_out_r_39__N_2714[1]), 
            .\pin_intrpt[7] (pin_intrpt[7])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(304[3] 325[2])
    cs_decoder u_cs_decoder (.cs_decoded({cs_decoded}), .CS_READY_c(CS_READY_c), 
            .FLASH_CS_c(FLASH_CS_c), .MAX3421_CS_c(MAX3421_CS_c), .cs_c_0(cs_c_0), 
            .cs_c_1(cs_c_1), .cs_c_2(cs_c_2), .cs_c_4(cs_c_4), .cs_c_3(cs_c_3)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(213[3] 221[2])
    \intrpt_ctrl(DEV_ID=1)  \intrpt_ins_1..u_intrpt_ctrl  (.clk(clk), .n29239(n29239), 
            .\spi_data_out_r_39__N_2643[0] (spi_data_out_r_39__N_2643[0]), 
            .\pin_intrpt[3] (pin_intrpt[3]), .intrpt_out_c_1(intrpt_out_c_1), 
            .intrpt_out_N_2706(intrpt_out_N_2706), .n29757(n29757), .clear_intrpt(clear_intrpt_adj_7956), 
            .clear_intrpt_N_2710(clear_intrpt_N_2710), .\spi_data_out_r_39__N_2643[2] (spi_data_out_r_39__N_2643[2]), 
            .\pin_intrpt[5] (pin_intrpt[5]), .\spi_data_out_r_39__N_2643[1] (spi_data_out_r_39__N_2643[1]), 
            .\pin_intrpt[4] (pin_intrpt[4])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(304[3] 325[2])
    intrpt_ctrl \intrpt_ins_0..u_intrpt_ctrl  (.\spi_data_out_r_39__N_2572[0] (spi_data_out_r_39__N_2572[0]), 
            .clk(clk), .\pin_intrpt[0] (pin_intrpt[0]), .n29239(n29239), 
            .intrpt_out_c_0(intrpt_out_c_0), .intrpt_out_N_2635(intrpt_out_N_2635), 
            .n29757(n29757), .clear_intrpt(clear_intrpt), .clear_intrpt_N_2639(clear_intrpt_N_2639), 
            .n29212(n29212), .\spi_cmd[2] (spi_cmd[2]), .n29126(n29126), 
            .\spi_addr[0] (spi_addr[0]), .clear_intrpt_N_2781(clear_intrpt_N_2781), 
            .clear_intrpt_N_2852(clear_intrpt_N_2852), .n29178(n29178), 
            .n29141(n29141), .\spi_cmd[1] (spi_cmd[1]), .clear_intrpt_N_2923(clear_intrpt_N_2923), 
            .clear_intrpt_N_2994(clear_intrpt_N_2994), .\spi_data_out_r_39__N_2572[2] (spi_data_out_r_39__N_2572[2]), 
            .\mode[2]_derived_32 (mode_2_derived_32), .\spi_data_out_r_39__N_2572[1] (spi_data_out_r_39__N_2572[1]), 
            .\pin_intrpt[1] (pin_intrpt[1]), .n29761(n29761), .\spi_addr[1] (spi_addr[1]), 
            .n29310(n29310), .\spi_addr[2] (spi_addr[2]), .n13413(n13413)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(304[3] 325[2])
    quad_decoder \quad_ins_0..u_quad_decoder  (.n29099(n29099), .n25293(n25293), 
            .quad_buffer({quad_buffer_adj_8522}), .quad_count({quad_count_adj_8521}), 
            .\spi_data_out_r_39__N_2483[9] (spi_data_out_r_39__N_2483[9]), 
            .\spi_data_out_r_39__N_2483[8] (spi_data_out_r_39__N_2483[8]), 
            .clk_1MHz(clk_1MHz), .clk_1MHz_enable_340(clk_1MHz_enable_340), 
            .\spi_data_out_r_39__N_934[0] (spi_data_out_r_39__N_934[0]), .clk(clk), 
            .\quad_b[0] (quad_b[0]), .\mode[2]_derived_32 (mode_2_derived_32), 
            .\spi_data_out_r_39__N_2483[7] (spi_data_out_r_39__N_2483[7]), 
            .\spi_data_out_r_39__N_2483[6] (spi_data_out_r_39__N_2483[6]), 
            .\spi_data_out_r_39__N_2483[5] (spi_data_out_r_39__N_2483[5]), 
            .\spi_data_out_r_39__N_2483[4] (spi_data_out_r_39__N_2483[4]), 
            .\spi_data_out_r_39__N_2483[3] (spi_data_out_r_39__N_2483[3]), 
            .\spi_data_out_r_39__N_2483[2] (spi_data_out_r_39__N_2483[2]), 
            .n13413(n13413), .quad_buffer_adj_528({quad_buffer_adj_8286}), 
            .quad_count_adj_529({quad_count_adj_8285}), .\spi_data_out_r_39__N_1547[29] (spi_data_out_r_39__N_1547[29]), 
            .\spi_data_out_r_39__N_2483[1] (spi_data_out_r_39__N_2483[1]), 
            .n29239(n29239), .\spi_addr[1] (spi_addr[1]), .n29761(n29761), 
            .\spi_addr[2] (spi_addr[2]), .n13506(n13506), .n13511(n13511), 
            .\spi_data_out_r_39__N_1547[28] (spi_data_out_r_39__N_1547[28]), 
            .clk_enable_433(clk_enable_433), .\spi_data_r[0] (spi_data_r[0]), 
            .quad_homing({quad_homing}), .clk_enable_436(clk_enable_436), 
            .n29762(n29762), .n29098(n29098), .quad_buffer_adj_530({quad_buffer_adj_8463}), 
            .quad_count_adj_531({quad_count_adj_8462}), .\spi_data_out_r_39__N_2249[0] (spi_data_out_r_39__N_2249[0]), 
            .\spi_data_out_r_39__N_2249[31] (spi_data_out_r_39__N_2249[31]), 
            .\spi_data_out_r_39__N_2249[30] (spi_data_out_r_39__N_2249[30]), 
            .\spi_data_out_r_39__N_2249[29] (spi_data_out_r_39__N_2249[29]), 
            .\spi_data_out_r_39__N_2249[28] (spi_data_out_r_39__N_2249[28]), 
            .\spi_data_out_r_39__N_2249[27] (spi_data_out_r_39__N_2249[27]), 
            .\spi_data_out_r_39__N_2249[26] (spi_data_out_r_39__N_2249[26]), 
            .\spi_data_out_r_39__N_2249[25] (spi_data_out_r_39__N_2249[25]), 
            .\spi_data_out_r_39__N_2249[24] (spi_data_out_r_39__N_2249[24]), 
            .\spi_data_out_r_39__N_2249[23] (spi_data_out_r_39__N_2249[23]), 
            .\spi_data_out_r_39__N_2249[22] (spi_data_out_r_39__N_2249[22]), 
            .\spi_data_out_r_39__N_1547[27] (spi_data_out_r_39__N_1547[27]), 
            .\spi_data_out_r_39__N_2249[21] (spi_data_out_r_39__N_2249[21]), 
            .\spi_data_out_r_39__N_2249[20] (spi_data_out_r_39__N_2249[20]), 
            .quad_buffer_adj_532({quad_buffer_adj_8404}), .quad_count_adj_533({quad_count_adj_8403}), 
            .\spi_data_out_r_39__N_2015[27] (spi_data_out_r_39__N_2015[27]), 
            .\spi_data_out_r_39__N_2015[26] (spi_data_out_r_39__N_2015[26]), 
            .\spi_data_out_r_39__N_2015[25] (spi_data_out_r_39__N_2015[25]), 
            .\spi_data_out_r_39__N_2015[24] (spi_data_out_r_39__N_2015[24]), 
            .\spi_data_out_r_39__N_2015[23] (spi_data_out_r_39__N_2015[23]), 
            .\spi_data_out_r_39__N_2249[19] (spi_data_out_r_39__N_2249[19]), 
            .\spi_data_out_r_39__N_2249[18] (spi_data_out_r_39__N_2249[18]), 
            .\spi_data_out_r_39__N_1547[26] (spi_data_out_r_39__N_1547[26]), 
            .\spi_data_out_r_39__N_1547[25] (spi_data_out_r_39__N_1547[25]), 
            .\spi_data_out_r_39__N_2249[17] (spi_data_out_r_39__N_2249[17]), 
            .\spi_data_out_r_39__N_2015[22] (spi_data_out_r_39__N_2015[22]), 
            .\spi_data_out_r_39__N_2249[16] (spi_data_out_r_39__N_2249[16]), 
            .\spi_data_out_r_39__N_2249[15] (spi_data_out_r_39__N_2249[15]), 
            .\spi_data_out_r_39__N_1547[24] (spi_data_out_r_39__N_1547[24]), 
            .\spi_data_out_r_39__N_2249[14] (spi_data_out_r_39__N_2249[14]), 
            .\spi_data_out_r_39__N_2015[21] (spi_data_out_r_39__N_2015[21]), 
            .\spi_data_out_r_39__N_2015[20] (spi_data_out_r_39__N_2015[20]), 
            .\spi_data_out_r_39__N_2249[13] (spi_data_out_r_39__N_2249[13]), 
            .\spi_data_out_r_39__N_2015[19] (spi_data_out_r_39__N_2015[19]), 
            .\spi_data_out_r_39__N_2015[18] (spi_data_out_r_39__N_2015[18]), 
            .\spi_data_out_r_39__N_2015[17] (spi_data_out_r_39__N_2015[17]), 
            .\spi_data_out_r_39__N_2249[12] (spi_data_out_r_39__N_2249[12]), 
            .\spi_data_out_r_39__N_2015[16] (spi_data_out_r_39__N_2015[16]), 
            .\spi_data_out_r_39__N_2015[15] (spi_data_out_r_39__N_2015[15]), 
            .\spi_data_out_r_39__N_2015[14] (spi_data_out_r_39__N_2015[14]), 
            .\spi_data_out_r_39__N_2015[13] (spi_data_out_r_39__N_2015[13]), 
            .\spi_data_out_r_39__N_2249[11] (spi_data_out_r_39__N_2249[11]), 
            .\spi_data_out_r_39__N_2249[10] (spi_data_out_r_39__N_2249[10]), 
            .\spi_data_out_r_39__N_2249[9] (spi_data_out_r_39__N_2249[9]), 
            .spi_data_out_r_39__N_974(spi_data_out_r_39__N_974), .spi_data_out_r_39__N_1162(spi_data_out_r_39__N_1162), 
            .\spi_data_out_r_39__N_2249[8] (spi_data_out_r_39__N_2249[8]), 
            .quad_set_complete(quad_set_complete), .quad_set_valid(quad_set_valid), 
            .\spi_data_out_r_39__N_2015[12] (spi_data_out_r_39__N_2015[12]), 
            .\spi_data_out_r_39__N_2015[11] (spi_data_out_r_39__N_2015[11]), 
            .\spi_data_out_r_39__N_2249[7] (spi_data_out_r_39__N_2249[7]), 
            .\spi_data_out_r_39__N_2249[6] (spi_data_out_r_39__N_2249[6]), 
            .\spi_data_out_r_39__N_2249[5] (spi_data_out_r_39__N_2249[5]), 
            .\spi_data_out_r_39__N_2249[4] (spi_data_out_r_39__N_2249[4]), 
            .\spi_data_out_r_39__N_1547[23] (spi_data_out_r_39__N_1547[23]), 
            .\spi_data_out_r_39__N_2015[10] (spi_data_out_r_39__N_2015[10]), 
            .\spi_data_out_r_39__N_2015[9] (spi_data_out_r_39__N_2015[9]), 
            .\spi_data_out_r_39__N_2249[3] (spi_data_out_r_39__N_2249[3]), 
            .\spi_data_out_r_39__N_2015[8] (spi_data_out_r_39__N_2015[8]), 
            .\spi_data_out_r_39__N_2015[7] (spi_data_out_r_39__N_2015[7]), 
            .\spi_data_out_r_39__N_2015[6] (spi_data_out_r_39__N_2015[6]), 
            .\spi_data_out_r_39__N_2015[5] (spi_data_out_r_39__N_2015[5]), 
            .\spi_data_out_r_39__N_1547[22] (spi_data_out_r_39__N_1547[22]), 
            .\spi_data_out_r_39__N_2249[2] (spi_data_out_r_39__N_2249[2]), 
            .\spi_data_out_r_39__N_1547[21] (spi_data_out_r_39__N_1547[21]), 
            .\spi_data_out_r_39__N_2015[4] (spi_data_out_r_39__N_2015[4]), 
            .\spi_data_out_r_39__N_2015[3] (spi_data_out_r_39__N_2015[3]), 
            .\spi_data_out_r_39__N_1547[20] (spi_data_out_r_39__N_1547[20]), 
            .\spi_data_out_r_39__N_2249[1] (spi_data_out_r_39__N_2249[1]), 
            .\spi_data_out_r_39__N_2015[2] (spi_data_out_r_39__N_2015[2]), 
            .\spi_data_out_r_39__N_2015[1] (spi_data_out_r_39__N_2015[1]), 
            .quad_buffer_adj_534({quad_buffer_adj_8345}), .quad_count_adj_535({quad_count_adj_8344}), 
            .\spi_data_out_r_39__N_1781[0] (spi_data_out_r_39__N_1781[0]), 
            .\spi_data_out_r_39__N_1547[19] (spi_data_out_r_39__N_1547[19]), 
            .\spi_data_out_r_39__N_1781[31] (spi_data_out_r_39__N_1781[31]), 
            .\spi_data_out_r_39__N_1781[30] (spi_data_out_r_39__N_1781[30]), 
            .\spi_data_out_r_39__N_1781[29] (spi_data_out_r_39__N_1781[29]), 
            .\spi_data_out_r_39__N_1781[28] (spi_data_out_r_39__N_1781[28]), 
            .\spi_data_out_r_39__N_1781[27] (spi_data_out_r_39__N_1781[27]), 
            .n29260(n29260), .pin_io_out_4(pin_io_out_4), .n108(n108), 
            .n79(n79), .\spi_data_out_r_39__N_1781[26] (spi_data_out_r_39__N_1781[26]), 
            .\spi_data_out_r_39__N_1547[18] (spi_data_out_r_39__N_1547[18]), 
            .\spi_data_out_r_39__N_1547[17] (spi_data_out_r_39__N_1547[17]), 
            .\spi_data_out_r_39__N_1781[25] (spi_data_out_r_39__N_1781[25]), 
            .\spi_data_out_r_39__N_1781[24] (spi_data_out_r_39__N_1781[24]), 
            .\spi_data_out_r_39__N_1781[23] (spi_data_out_r_39__N_1781[23]), 
            .\spi_data_out_r_39__N_1547[16] (spi_data_out_r_39__N_1547[16]), 
            .\spi_data_out_r_39__N_1781[22] (spi_data_out_r_39__N_1781[22]), 
            .\spi_data_out_r_39__N_1781[21] (spi_data_out_r_39__N_1781[21]), 
            .\spi_data_out_r_39__N_1781[20] (spi_data_out_r_39__N_1781[20]), 
            .\spi_data_out_r_39__N_1781[19] (spi_data_out_r_39__N_1781[19]), 
            .\spi_data_out_r_39__N_1781[18] (spi_data_out_r_39__N_1781[18]), 
            .\spi_data_out_r_39__N_1547[15] (spi_data_out_r_39__N_1547[15]), 
            .\spi_data_out_r_39__N_1547[14] (spi_data_out_r_39__N_1547[14]), 
            .\spi_data_out_r_39__N_1781[17] (spi_data_out_r_39__N_1781[17]), 
            .\spi_data_out_r_39__N_1781[16] (spi_data_out_r_39__N_1781[16]), 
            .\spi_data_out_r_39__N_1781[15] (spi_data_out_r_39__N_1781[15]), 
            .\spi_data_out_r_39__N_1781[14] (spi_data_out_r_39__N_1781[14]), 
            .\spi_data_out_r_39__N_1781[13] (spi_data_out_r_39__N_1781[13]), 
            .\spi_data_out_r_39__N_1781[12] (spi_data_out_r_39__N_1781[12]), 
            .\spi_data_out_r_39__N_1781[11] (spi_data_out_r_39__N_1781[11]), 
            .\spi_data_out_r_39__N_1547[13] (spi_data_out_r_39__N_1547[13]), 
            .\spi_data_out_r_39__N_1781[10] (spi_data_out_r_39__N_1781[10]), 
            .\spi_data_out_r_39__N_1781[9] (spi_data_out_r_39__N_1781[9]), 
            .\spi_data_out_r_39__N_1781[8] (spi_data_out_r_39__N_1781[8]), 
            .\spi_data_out_r_39__N_1781[7] (spi_data_out_r_39__N_1781[7]), 
            .\spi_data_out_r_39__N_1781[6] (spi_data_out_r_39__N_1781[6]), 
            .\spi_data_out_r_39__N_1781[5] (spi_data_out_r_39__N_1781[5]), 
            .n27256(n27256), .n29078(n29078), .n27338(n27338), .n29213(n29213), 
            .clk_enable_199(clk_enable_199), .\spi_data_out_r_39__N_1781[4] (spi_data_out_r_39__N_1781[4]), 
            .\spi_data_out_r_39__N_1781[3] (spi_data_out_r_39__N_1781[3]), 
            .\spi_data_out_r_39__N_1781[2] (spi_data_out_r_39__N_1781[2]), 
            .\spi_data_out_r_39__N_1781[1] (spi_data_out_r_39__N_1781[1]), 
            .\spi_data_out_r_39__N_2483[0] (spi_data_out_r_39__N_2483[0]), 
            .\spi_data_out_r_39__N_2483[31] (spi_data_out_r_39__N_2483[31]), 
            .\spi_data_out_r_39__N_2483[30] (spi_data_out_r_39__N_2483[30]), 
            .\spi_data_out_r_39__N_2483[29] (spi_data_out_r_39__N_2483[29]), 
            .\spi_data_out_r_39__N_2483[28] (spi_data_out_r_39__N_2483[28]), 
            .\spi_data_out_r_39__N_1547[0] (spi_data_out_r_39__N_1547[0]), 
            .\spi_data_out_r_39__N_2483[27] (spi_data_out_r_39__N_2483[27]), 
            .\spi_data_out_r_39__N_2483[26] (spi_data_out_r_39__N_2483[26]), 
            .resetn_c(resetn_c), .GND_net(GND_net), .\spi_data_out_r_39__N_2483[25] (spi_data_out_r_39__N_2483[25]), 
            .\spi_data_out_r_39__N_2483[24] (spi_data_out_r_39__N_2483[24]), 
            .\spi_data_out_r_39__N_2483[23] (spi_data_out_r_39__N_2483[23]), 
            .\spi_data_out_r_39__N_2483[22] (spi_data_out_r_39__N_2483[22]), 
            .\spi_data_out_r_39__N_2483[21] (spi_data_out_r_39__N_2483[21]), 
            .\spi_data_out_r_39__N_2483[20] (spi_data_out_r_39__N_2483[20]), 
            .\spi_data_out_r_39__N_2483[19] (spi_data_out_r_39__N_2483[19]), 
            .\spi_data_out_r_39__N_2483[18] (spi_data_out_r_39__N_2483[18]), 
            .\spi_data_out_r_39__N_2483[17] (spi_data_out_r_39__N_2483[17]), 
            .\spi_data_out_r_39__N_1547[12] (spi_data_out_r_39__N_1547[12]), 
            .\spi_data_out_r_39__N_2483[16] (spi_data_out_r_39__N_2483[16]), 
            .\spi_data_out_r_39__N_1547[31] (spi_data_out_r_39__N_1547[31]), 
            .\spi_data_out_r_39__N_2483[15] (spi_data_out_r_39__N_2483[15]), 
            .\spi_data_out_r_39__N_1547[30] (spi_data_out_r_39__N_1547[30]), 
            .\spi_data_out_r_39__N_2483[14] (spi_data_out_r_39__N_2483[14]), 
            .\spi_data_out_r_39__N_1547[11] (spi_data_out_r_39__N_1547[11]), 
            .\spi_data_out_r_39__N_1547[10] (spi_data_out_r_39__N_1547[10]), 
            .\spi_data_out_r_39__N_2483[13] (spi_data_out_r_39__N_2483[13]), 
            .\spi_data_out_r_39__N_1547[9] (spi_data_out_r_39__N_1547[9]), 
            .\spi_data_out_r_39__N_2483[12] (spi_data_out_r_39__N_2483[12]), 
            .\spi_data_out_r_39__N_2483[11] (spi_data_out_r_39__N_2483[11]), 
            .\spi_data_out_r_39__N_2483[10] (spi_data_out_r_39__N_2483[10]), 
            .\spi_data_out_r_39__N_1547[8] (spi_data_out_r_39__N_1547[8]), 
            .\quad_a[0] (quad_a[0]), .\spi_data_out_r_39__N_934[31] (spi_data_out_r_39__N_934[31]), 
            .\spi_data_out_r_39__N_934[30] (spi_data_out_r_39__N_934[30]), 
            .\spi_data_out_r_39__N_934[29] (spi_data_out_r_39__N_934[29]), 
            .\spi_data_out_r_39__N_1547[7] (spi_data_out_r_39__N_1547[7]), 
            .\spi_data_out_r_39__N_934[28] (spi_data_out_r_39__N_934[28]), 
            .\spi_data_out_r_39__N_934[27] (spi_data_out_r_39__N_934[27]), 
            .\spi_data_out_r_39__N_934[26] (spi_data_out_r_39__N_934[26]), 
            .\spi_data_out_r_39__N_934[25] (spi_data_out_r_39__N_934[25]), 
            .\spi_data_out_r_39__N_934[24] (spi_data_out_r_39__N_934[24]), 
            .\spi_data_out_r_39__N_934[23] (spi_data_out_r_39__N_934[23]), 
            .\spi_data_out_r_39__N_934[22] (spi_data_out_r_39__N_934[22]), 
            .\spi_data_out_r_39__N_934[21] (spi_data_out_r_39__N_934[21]), 
            .\spi_data_out_r_39__N_934[20] (spi_data_out_r_39__N_934[20]), 
            .\spi_data_out_r_39__N_934[19] (spi_data_out_r_39__N_934[19]), 
            .\spi_data_out_r_39__N_934[18] (spi_data_out_r_39__N_934[18]), 
            .\spi_data_out_r_39__N_934[17] (spi_data_out_r_39__N_934[17]), 
            .\spi_data_out_r_39__N_934[16] (spi_data_out_r_39__N_934[16]), 
            .\spi_data_out_r_39__N_934[15] (spi_data_out_r_39__N_934[15]), 
            .\spi_data_out_r_39__N_934[14] (spi_data_out_r_39__N_934[14]), 
            .\spi_data_out_r_39__N_934[13] (spi_data_out_r_39__N_934[13]), 
            .\spi_data_out_r_39__N_934[12] (spi_data_out_r_39__N_934[12]), 
            .\spi_data_out_r_39__N_934[11] (spi_data_out_r_39__N_934[11]), 
            .\spi_data_out_r_39__N_934[10] (spi_data_out_r_39__N_934[10]), 
            .\spi_data_out_r_39__N_934[9] (spi_data_out_r_39__N_934[9]), .\spi_data_out_r_39__N_934[8] (spi_data_out_r_39__N_934[8]), 
            .\spi_data_out_r_39__N_934[7] (spi_data_out_r_39__N_934[7]), .\spi_data_out_r_39__N_934[6] (spi_data_out_r_39__N_934[6]), 
            .\spi_data_out_r_39__N_934[5] (spi_data_out_r_39__N_934[5]), .\spi_data_out_r_39__N_934[4] (spi_data_out_r_39__N_934[4]), 
            .\spi_data_out_r_39__N_934[3] (spi_data_out_r_39__N_934[3]), .\spi_data_out_r_39__N_934[2] (spi_data_out_r_39__N_934[2]), 
            .\spi_data_out_r_39__N_934[1] (spi_data_out_r_39__N_934[1]), .\spi_data_out_r_39__N_1547[6] (spi_data_out_r_39__N_1547[6]), 
            .\spi_data_out_r_39__N_1547[5] (spi_data_out_r_39__N_1547[5]), 
            .\spi_data_out_r_39__N_1547[4] (spi_data_out_r_39__N_1547[4]), 
            .\spi_data_out_r_39__N_1547[3] (spi_data_out_r_39__N_1547[3]), 
            .\spi_data_out_r_39__N_1547[2] (spi_data_out_r_39__N_1547[2]), 
            .\spi_data_out_r_39__N_1547[1] (spi_data_out_r_39__N_1547[1]), 
            .quad_buffer_adj_536({quad_buffer_adj_8227}), .quad_count_adj_537({quad_count_adj_8226}), 
            .\spi_data_out_r_39__N_1313[0] (spi_data_out_r_39__N_1313[0]), 
            .\spi_data_out_r_39__N_1313[31] (spi_data_out_r_39__N_1313[31]), 
            .\spi_cmd[2] (spi_cmd[2]), .n29117(n29117), .n29310(n29310), 
            .clear_intrpt_N_3065(clear_intrpt_N_3065), .\spi_data_out_r_39__N_1313[30] (spi_data_out_r_39__N_1313[30]), 
            .\spi_data_out_r_39__N_1313[29] (spi_data_out_r_39__N_1313[29]), 
            .\spi_data_out_r_39__N_1313[28] (spi_data_out_r_39__N_1313[28]), 
            .\spi_data_out_r_39__N_1313[27] (spi_data_out_r_39__N_1313[27]), 
            .\spi_data_r[1] (spi_data_r[1]), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[3] (spi_data_r[3]), .\spi_data_r[4] (spi_data_r[4]), 
            .\spi_data_r[5] (spi_data_r[5]), .\spi_data_r[6] (spi_data_r[6]), 
            .\spi_data_r[7] (spi_data_r[7]), .\spi_data_r[8] (spi_data_r[8]), 
            .\spi_data_r[9] (spi_data_r[9]), .\spi_data_r[10] (spi_data_r[10]), 
            .\spi_data_r[11] (spi_data_r[11]), .\spi_data_r[12] (spi_data_r[12]), 
            .\spi_data_r[13] (spi_data_r[13]), .\spi_data_r[14] (spi_data_r[14]), 
            .\spi_data_r[15] (spi_data_r[15]), .\spi_data_r[16] (spi_data_r[16]), 
            .\spi_data_r[17] (spi_data_r[17]), .\spi_data_r[18] (spi_data_r[18]), 
            .\spi_data_r[19] (spi_data_r[19]), .\spi_data_r[20] (spi_data_r[20]), 
            .\spi_data_r[21] (spi_data_r[21]), .\spi_data_r[22] (spi_data_r[22]), 
            .\spi_data_r[23] (spi_data_r[23]), .\spi_data_r[24] (spi_data_r[24]), 
            .\spi_data_r[25] (spi_data_r[25]), .\spi_data_r[26] (spi_data_r[26]), 
            .\spi_data_r[27] (spi_data_r[27]), .\spi_data_r[28] (spi_data_r[28]), 
            .\spi_data_r[29] (spi_data_r[29]), .\spi_data_r[30] (spi_data_r[30]), 
            .\spi_data_r[31] (spi_data_r[31]), .clk_enable_501(clk_enable_501), 
            .n29085(n29085), .\spi_data_out_r_39__N_1313[26] (spi_data_out_r_39__N_1313[26]), 
            .\spi_data_out_r_39__N_1313[25] (spi_data_out_r_39__N_1313[25]), 
            .\spi_data_out_r_39__N_1313[24] (spi_data_out_r_39__N_1313[24]), 
            .n3(n3), .n26(n26), .\spi_data_out_r_39__N_1313[23] (spi_data_out_r_39__N_1313[23]), 
            .\spi_data_out_r_39__N_1313[22] (spi_data_out_r_39__N_1313[22]), 
            .\spi_data_out_r_39__N_1313[21] (spi_data_out_r_39__N_1313[21]), 
            .\spi_data_out_r_39__N_1313[20] (spi_data_out_r_39__N_1313[20]), 
            .\spi_data_out_r_39__N_1313[19] (spi_data_out_r_39__N_1313[19]), 
            .\spi_data_out_r_39__N_1313[18] (spi_data_out_r_39__N_1313[18]), 
            .\spi_data_out_r_39__N_1313[17] (spi_data_out_r_39__N_1313[17]), 
            .n20819(n20819), .\spi_data_out_r_39__N_1313[16] (spi_data_out_r_39__N_1313[16]), 
            .\spi_data_out_r_39__N_1313[15] (spi_data_out_r_39__N_1313[15]), 
            .\spi_data_out_r_39__N_1313[14] (spi_data_out_r_39__N_1313[14]), 
            .n31(n31), .\spi_data_out_r_39__N_1313[13] (spi_data_out_r_39__N_1313[13]), 
            .\spi_data_out_r_39__N_1313[12] (spi_data_out_r_39__N_1313[12]), 
            .\spi_data_out_r_39__N_1313[11] (spi_data_out_r_39__N_1313[11]), 
            .\spi_data_out_r_39__N_1313[10] (spi_data_out_r_39__N_1313[10]), 
            .\spi_data_out_r_39__N_1313[9] (spi_data_out_r_39__N_1313[9]), 
            .\spi_data_out_r_39__N_1313[8] (spi_data_out_r_39__N_1313[8]), 
            .\spi_data_out_r_39__N_1313[7] (spi_data_out_r_39__N_1313[7]), 
            .\spi_data_out_r_39__N_1313[6] (spi_data_out_r_39__N_1313[6]), 
            .\spi_data_out_r_39__N_1313[5] (spi_data_out_r_39__N_1313[5]), 
            .\spi_data_out_r_39__N_1313[4] (spi_data_out_r_39__N_1313[4]), 
            .\spi_data_out_r_39__N_1313[3] (spi_data_out_r_39__N_1313[3]), 
            .\spi_data_out_r_39__N_1313[2] (spi_data_out_r_39__N_1313[2]), 
            .\spi_data_out_r_39__N_1313[1] (spi_data_out_r_39__N_1313[1]), 
            .\spi_data_out_r_39__N_2015[0] (spi_data_out_r_39__N_2015[0]), 
            .\spi_data_out_r_39__N_2015[31] (spi_data_out_r_39__N_2015[31]), 
            .\spi_data_out_r_39__N_2015[30] (spi_data_out_r_39__N_2015[30]), 
            .\spi_data_out_r_39__N_2015[29] (spi_data_out_r_39__N_2015[29]), 
            .n29326(n29326), .\spi_data_out_r_39__N_2015[28] (spi_data_out_r_39__N_2015[28])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(272[3] 293[2])
    \quad_decoder(DEV_ID=2)  \quad_ins_2..u_quad_decoder  (.quad_count({quad_count_adj_8285}), 
            .clk_1MHz(clk_1MHz), .\spi_data_out_r_39__N_1402[0] (spi_data_out_r_39__N_1402[0]), 
            .clk(clk), .\spi_data_out_r_39__N_1547[0] (spi_data_out_r_39__N_1547[0]), 
            .\quad_b[2] (quad_b[2]), .quad_buffer({quad_buffer_adj_8286}), 
            .\mode[2]_derived_32 (mode_2_derived_32_adj_8013), .clk_enable_269(clk_enable_269), 
            .n29239(n29239), .\spi_data_r[0] (spi_data_r[0]), .n26948(n26948), 
            .quad_homing({quad_homing_adj_8284}), .clk_enable_435(clk_enable_435), 
            .n29762(n29762), .spi_data_out_r_39__N_1442(spi_data_out_r_39__N_1442), 
            .quad_set_complete(quad_set_complete_adj_7623), .n29099(n29099), 
            .\spi_addr[0] (spi_addr[0]), .n26933(n26933), .n13506(n13506), 
            .spi_data_out_r_39__N_1162(spi_data_out_r_39__N_1162), .n13413(n13413), 
            .resetn_c(resetn_c), .n13511(n13511), .spi_data_out_r_39__N_2098(spi_data_out_r_39__N_2098), 
            .n25293(n25293), .spi_data_out_r_39__N_2566(spi_data_out_r_39__N_2566), 
            .pin_io_out_24(pin_io_out_24), .n29233(n29233), .\spi_data_r[31] (spi_data_r[31]), 
            .\spi_data_r[30] (spi_data_r[30]), .\spi_data_r[29] (spi_data_r[29]), 
            .\spi_data_r[28] (spi_data_r[28]), .\spi_data_r[27] (spi_data_r[27]), 
            .\spi_data_r[26] (spi_data_r[26]), .\spi_data_r[25] (spi_data_r[25]), 
            .\spi_data_r[24] (spi_data_r[24]), .\spi_data_r[23] (spi_data_r[23]), 
            .\spi_data_r[22] (spi_data_r[22]), .\spi_data_r[21] (spi_data_r[21]), 
            .\spi_data_r[20] (spi_data_r[20]), .\spi_data_r[19] (spi_data_r[19]), 
            .\spi_data_r[18] (spi_data_r[18]), .\spi_data_r[17] (spi_data_r[17]), 
            .\spi_data_r[16] (spi_data_r[16]), .\spi_data_r[15] (spi_data_r[15]), 
            .\spi_data_r[14] (spi_data_r[14]), .\spi_data_r[13] (spi_data_r[13]), 
            .\spi_data_r[12] (spi_data_r[12]), .\spi_data_r[11] (spi_data_r[11]), 
            .\spi_data_r[10] (spi_data_r[10]), .\spi_data_r[9] (spi_data_r[9]), 
            .\spi_data_r[8] (spi_data_r[8]), .\spi_data_r[7] (spi_data_r[7]), 
            .\spi_data_r[6] (spi_data_r[6]), .\spi_data_r[5] (spi_data_r[5]), 
            .\spi_data_r[4] (spi_data_r[4]), .\spi_data_r[3] (spi_data_r[3]), 
            .\spi_data_r[2] (spi_data_r[2]), .\spi_data_r[1] (spi_data_r[1]), 
            .\quad_a[2] (quad_a[2]), .\spi_data_out_r_39__N_1402[31] (spi_data_out_r_39__N_1402[31]), 
            .\spi_data_out_r_39__N_1547[31] (spi_data_out_r_39__N_1547[31]), 
            .\spi_data_out_r_39__N_1402[30] (spi_data_out_r_39__N_1402[30]), 
            .\spi_data_out_r_39__N_1547[30] (spi_data_out_r_39__N_1547[30]), 
            .\spi_data_out_r_39__N_1402[29] (spi_data_out_r_39__N_1402[29]), 
            .\spi_data_out_r_39__N_1547[29] (spi_data_out_r_39__N_1547[29]), 
            .\spi_data_out_r_39__N_1402[28] (spi_data_out_r_39__N_1402[28]), 
            .\spi_data_out_r_39__N_1547[28] (spi_data_out_r_39__N_1547[28]), 
            .\spi_data_out_r_39__N_1402[27] (spi_data_out_r_39__N_1402[27]), 
            .\spi_data_out_r_39__N_1547[27] (spi_data_out_r_39__N_1547[27]), 
            .\spi_data_out_r_39__N_1402[26] (spi_data_out_r_39__N_1402[26]), 
            .\spi_data_out_r_39__N_1547[26] (spi_data_out_r_39__N_1547[26]), 
            .\spi_data_out_r_39__N_1402[25] (spi_data_out_r_39__N_1402[25]), 
            .\spi_data_out_r_39__N_1547[25] (spi_data_out_r_39__N_1547[25]), 
            .\spi_data_out_r_39__N_1402[24] (spi_data_out_r_39__N_1402[24]), 
            .\spi_data_out_r_39__N_1547[24] (spi_data_out_r_39__N_1547[24]), 
            .\spi_data_out_r_39__N_1402[23] (spi_data_out_r_39__N_1402[23]), 
            .\spi_data_out_r_39__N_1547[23] (spi_data_out_r_39__N_1547[23]), 
            .\spi_data_out_r_39__N_1402[22] (spi_data_out_r_39__N_1402[22]), 
            .\spi_data_out_r_39__N_1547[22] (spi_data_out_r_39__N_1547[22]), 
            .\spi_data_out_r_39__N_1402[21] (spi_data_out_r_39__N_1402[21]), 
            .\spi_data_out_r_39__N_1547[21] (spi_data_out_r_39__N_1547[21]), 
            .\spi_data_out_r_39__N_1402[20] (spi_data_out_r_39__N_1402[20]), 
            .\spi_data_out_r_39__N_1547[20] (spi_data_out_r_39__N_1547[20]), 
            .\spi_data_out_r_39__N_1402[19] (spi_data_out_r_39__N_1402[19]), 
            .\spi_data_out_r_39__N_1547[19] (spi_data_out_r_39__N_1547[19]), 
            .\spi_data_out_r_39__N_1402[18] (spi_data_out_r_39__N_1402[18]), 
            .\spi_data_out_r_39__N_1547[18] (spi_data_out_r_39__N_1547[18]), 
            .\spi_data_out_r_39__N_1402[17] (spi_data_out_r_39__N_1402[17]), 
            .\spi_data_out_r_39__N_1547[17] (spi_data_out_r_39__N_1547[17]), 
            .\spi_data_out_r_39__N_1402[16] (spi_data_out_r_39__N_1402[16]), 
            .\spi_data_out_r_39__N_1547[16] (spi_data_out_r_39__N_1547[16]), 
            .\spi_data_out_r_39__N_1402[15] (spi_data_out_r_39__N_1402[15]), 
            .\spi_data_out_r_39__N_1547[15] (spi_data_out_r_39__N_1547[15]), 
            .\spi_data_out_r_39__N_1402[14] (spi_data_out_r_39__N_1402[14]), 
            .\spi_data_out_r_39__N_1547[14] (spi_data_out_r_39__N_1547[14]), 
            .\spi_data_out_r_39__N_1402[13] (spi_data_out_r_39__N_1402[13]), 
            .\spi_data_out_r_39__N_1547[13] (spi_data_out_r_39__N_1547[13]), 
            .\spi_data_out_r_39__N_1402[12] (spi_data_out_r_39__N_1402[12]), 
            .\spi_data_out_r_39__N_1547[12] (spi_data_out_r_39__N_1547[12]), 
            .\spi_data_out_r_39__N_1402[11] (spi_data_out_r_39__N_1402[11]), 
            .\spi_data_out_r_39__N_1547[11] (spi_data_out_r_39__N_1547[11]), 
            .\spi_data_out_r_39__N_1402[10] (spi_data_out_r_39__N_1402[10]), 
            .\spi_data_out_r_39__N_1547[10] (spi_data_out_r_39__N_1547[10]), 
            .\spi_data_out_r_39__N_1402[9] (spi_data_out_r_39__N_1402[9]), 
            .\spi_data_out_r_39__N_1547[9] (spi_data_out_r_39__N_1547[9]), 
            .\spi_data_out_r_39__N_1402[8] (spi_data_out_r_39__N_1402[8]), 
            .\spi_data_out_r_39__N_1547[8] (spi_data_out_r_39__N_1547[8]), 
            .\spi_data_out_r_39__N_1402[7] (spi_data_out_r_39__N_1402[7]), 
            .\spi_data_out_r_39__N_1547[7] (spi_data_out_r_39__N_1547[7]), 
            .\spi_data_out_r_39__N_1402[6] (spi_data_out_r_39__N_1402[6]), 
            .\spi_data_out_r_39__N_1547[6] (spi_data_out_r_39__N_1547[6]), 
            .\spi_data_out_r_39__N_1402[5] (spi_data_out_r_39__N_1402[5]), 
            .\spi_data_out_r_39__N_1547[5] (spi_data_out_r_39__N_1547[5]), 
            .\spi_data_out_r_39__N_1402[4] (spi_data_out_r_39__N_1402[4]), 
            .\spi_data_out_r_39__N_1547[4] (spi_data_out_r_39__N_1547[4]), 
            .\spi_data_out_r_39__N_1402[3] (spi_data_out_r_39__N_1402[3]), 
            .\spi_data_out_r_39__N_1547[3] (spi_data_out_r_39__N_1547[3]), 
            .\spi_data_out_r_39__N_1402[2] (spi_data_out_r_39__N_1402[2]), 
            .\spi_data_out_r_39__N_1547[2] (spi_data_out_r_39__N_1547[2]), 
            .\spi_data_out_r_39__N_1402[1] (spi_data_out_r_39__N_1402[1]), 
            .\spi_data_out_r_39__N_1547[1] (spi_data_out_r_39__N_1547[1]), 
            .n27301(n27301), .clk_enable_503(clk_enable_503), .n29122(n29122), 
            .GND_net(GND_net), .n29326(n29326), .n108(n108), .quad_set_valid(quad_set_valid), 
            .n3(n3), .mem_rdata_update_N_729(mem_rdata_update_N_729), .n9633(n9633), 
            .n12714(n12714), .n13(n13_adj_7890), .n29336(n29336), .n95(n95), 
            .quad_set_valid_adj_207(quad_set_valid_adj_7824), .n5647(n5647)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(272[3] 293[2])
    pll __ (.clk_in_c(clk_in_c), .clk_1MHz(clk_1MHz), .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(149[5:100])
    LUT4 i22830_2_lut (.A(n19361), .B(resetn_c), .Z(clk_1MHz_enable_24)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i22830_2_lut.init = 16'h7777;
    \piezo(DEV_ID=6,UART_ADDRESS_WIDTH=4)  \piezo_ins_6..u_piezo  (.n28811(n28811), 
            .n28813(n28813), .mode(mode_adj_8150), .clk(clk), .clk_enable_188(clk_enable_188), 
            .n29239(n29239), .n29762(n29762), .n29191(n29191), .n29190(n29190), 
            .pin_io_out_65(pin_io_out_65), .n25382(n25382), .pin_io_out_26(pin_io_out_26), 
            .pin_io_out_16(pin_io_out_16), .n29157(n29157), .n7(n7), .pin_io_out_40(pin_io_out_40), 
            .n29189(n29189), .C_8_c(C_8_c), .tx_N_6443(tx_N_6443), .pin_io_out_45(pin_io_out_45), 
            .n27189(n27189), .pin_io_out_46(pin_io_out_46), .pin_io_out_55(pin_io_out_55), 
            .n29150(n29150), .n27186(n27186), .n29202(n29202), .pin_io_out_15(pin_io_out_15), 
            .n29198(n29198), .n13(n13_adj_8151), .pin_io_out_56(pin_io_out_56), 
            .n29196(n29196), .n29158(n29158), .n26972(n26972), .n22(n22), 
            .pin_io_out_5(pin_io_out_5), .n29160(n29160), .n29153(n29153), 
            .n26951(n26951), .n14(n14), .OW_ID_N_4464(OW_ID_N_4464), .n27480(n27480), 
            .n27483(n27483), .n29132(n29132), .n27471(n27471), .n29199(n29199), 
            .n27477(n27477), .mode_adj_183(mode_adj_8141), .mode_adj_184(mode_adj_8139), 
            .n29203(n29203), .mode_adj_185(mode_adj_8147), .mode_adj_186(mode_adj_8131), 
            .C_2_c_1(C_2_c_1), .C_1_c_0(C_1_c_0), .C_5_c_c(C_5_c_c), .n29313(n29313), 
            .mode_adj_187(mode_adj_8123), .n29284(n29284), .mode_adj_188(mode_adj_8137), 
            .mode_adj_189(mode_adj_8129), .mode_adj_190(mode_adj_8145), 
            .pin_io_out_25(pin_io_out_25), .n22_adj_191(n22_adj_7754), .mode_adj_192(mode_adj_8135), 
            .mode_adj_193(mode_adj_8144), .n31(n31_adj_8085), .mode_adj_194(mode_adj_8148), 
            .mode_adj_195(mode_adj_8132), .n29285(n29285), .\cs_decoded[8] (cs_decoded[8]), 
            .n5(n5), .mode_adj_196(mode_adj_8134), .n29293(n29293), .mode_adj_197(mode_adj_8149), 
            .mode_adj_198(mode_adj_8133), .n29299(n29299), .n29301(n29301), 
            .\mode[0] (n29785[0]), .n8679(n8679), .n29305(n29305), .\mode[1] (n29785[1]), 
            .n29300(n29300), .n29317(n29317), .n8739(n8739), .\cs_decoded[6] (cs_decoded[6]), 
            .n8740(n8740), .mode_adj_199(mode_adj_8130), .mode_adj_200(mode_adj_8146), 
            .n29303(n29303), .\cs_decoded[4] (cs_decoded[4]), .n29295(n29295), 
            .n8768(n8768), .\cs_decoded[13] (cs_decoded[13]), .n2(n2_adj_8155), 
            .n8836(n8836), .mode_adj_206({n29786}), .digital_output_r(digital_output_r_adj_8090), 
            .n26521(n26521), .n29267(n29267), .mode_adj_203(mode_adj_8142), 
            .pin_io_out_66(pin_io_out_66), .mode_adj_204(mode_adj_8127), 
            .pin_io_out_36(pin_io_out_36), .mode_adj_205(mode_adj_8124)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(632[3] 661[2])
    \intrpt_ctrl(DEV_ID=6)  \intrpt_ins_6..u_intrpt_ctrl  (.clk(clk), .n29239(n29239), 
            .\spi_data_out_r_39__N_2998[0] (spi_data_out_r_39__N_2998[0]), 
            .\pin_intrpt[18] (pin_intrpt[18]), .\pin_intrpt[20] (pin_intrpt[20]), 
            .\pin_intrpt[19] (pin_intrpt[19]), .clear_intrpt(clear_intrpt_adj_7962), 
            .clear_intrpt_N_3065(clear_intrpt_N_3065), .intrpt_out_c_6(intrpt_out_c_6), 
            .intrpt_out_N_3061(intrpt_out_N_3061), .n29757(n29757), .\spi_data_out_r_39__N_2998[2] (spi_data_out_r_39__N_2998[2]), 
            .\spi_data_out_r_39__N_2998[1] (spi_data_out_r_39__N_2998[1])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(304[3] 325[2])
    \quad_decoder(DEV_ID=3)  \quad_ins_3..u_quad_decoder  (.quad_count({quad_count_adj_8344}), 
            .clk_1MHz(clk_1MHz), .\spi_data_out_r_39__N_1636[0] (spi_data_out_r_39__N_1636[0]), 
            .clk(clk), .\spi_data_out_r_39__N_1781[0] (spi_data_out_r_39__N_1781[0]), 
            .\quad_b[3] (quad_b[3]), .quad_buffer({quad_buffer_adj_8345}), 
            .\pin_intrpt[11] (pin_intrpt[11]), .clk_enable_398(clk_enable_398), 
            .n29239(n29239), .\spi_data_r[0] (spi_data_r[0]), .clk_enable_434(clk_enable_434), 
            .n29762(n29762), .quad_set_complete(quad_set_complete_adj_7689), 
            .spi_data_out_r_39__N_1676(spi_data_out_r_39__N_1676), .n29098(n29098), 
            .\spi_addr[0] (spi_addr[0]), .n26933(n26933), .n13511(n13511), 
            .spi_data_out_r_39__N_2332(spi_data_out_r_39__N_2332), .n13506(n13506), 
            .spi_data_out_r_39__N_1396(spi_data_out_r_39__N_1396), .n13413(n13413), 
            .\quad_a[3] (quad_a[3]), .\spi_data_out_r_39__N_1636[31] (spi_data_out_r_39__N_1636[31]), 
            .\spi_data_out_r_39__N_1781[31] (spi_data_out_r_39__N_1781[31]), 
            .resetn_c(resetn_c), .GND_net(GND_net), .\spi_data_out_r_39__N_1636[30] (spi_data_out_r_39__N_1636[30]), 
            .\spi_data_out_r_39__N_1781[30] (spi_data_out_r_39__N_1781[30]), 
            .\spi_data_out_r_39__N_1636[29] (spi_data_out_r_39__N_1636[29]), 
            .\spi_data_out_r_39__N_1781[29] (spi_data_out_r_39__N_1781[29]), 
            .\spi_data_out_r_39__N_1636[28] (spi_data_out_r_39__N_1636[28]), 
            .\spi_data_out_r_39__N_1781[28] (spi_data_out_r_39__N_1781[28]), 
            .\spi_data_out_r_39__N_1636[27] (spi_data_out_r_39__N_1636[27]), 
            .\spi_data_out_r_39__N_1781[27] (spi_data_out_r_39__N_1781[27]), 
            .\spi_data_out_r_39__N_1636[26] (spi_data_out_r_39__N_1636[26]), 
            .\spi_data_out_r_39__N_1781[26] (spi_data_out_r_39__N_1781[26]), 
            .\spi_data_out_r_39__N_1636[25] (spi_data_out_r_39__N_1636[25]), 
            .\spi_data_out_r_39__N_1781[25] (spi_data_out_r_39__N_1781[25]), 
            .\spi_data_out_r_39__N_1636[24] (spi_data_out_r_39__N_1636[24]), 
            .\spi_data_out_r_39__N_1781[24] (spi_data_out_r_39__N_1781[24]), 
            .\spi_data_out_r_39__N_1636[23] (spi_data_out_r_39__N_1636[23]), 
            .\spi_data_out_r_39__N_1781[23] (spi_data_out_r_39__N_1781[23]), 
            .\spi_data_out_r_39__N_1636[22] (spi_data_out_r_39__N_1636[22]), 
            .\spi_data_out_r_39__N_1781[22] (spi_data_out_r_39__N_1781[22]), 
            .\spi_data_out_r_39__N_1636[21] (spi_data_out_r_39__N_1636[21]), 
            .\spi_data_out_r_39__N_1781[21] (spi_data_out_r_39__N_1781[21]), 
            .\spi_data_out_r_39__N_1636[20] (spi_data_out_r_39__N_1636[20]), 
            .\spi_data_out_r_39__N_1781[20] (spi_data_out_r_39__N_1781[20]), 
            .\spi_data_out_r_39__N_1636[19] (spi_data_out_r_39__N_1636[19]), 
            .\spi_data_out_r_39__N_1781[19] (spi_data_out_r_39__N_1781[19]), 
            .\spi_data_out_r_39__N_1636[18] (spi_data_out_r_39__N_1636[18]), 
            .\spi_data_out_r_39__N_1781[18] (spi_data_out_r_39__N_1781[18]), 
            .\spi_data_out_r_39__N_1636[17] (spi_data_out_r_39__N_1636[17]), 
            .\spi_data_out_r_39__N_1781[17] (spi_data_out_r_39__N_1781[17]), 
            .\spi_data_out_r_39__N_1636[16] (spi_data_out_r_39__N_1636[16]), 
            .\spi_data_out_r_39__N_1781[16] (spi_data_out_r_39__N_1781[16]), 
            .\spi_data_out_r_39__N_1636[15] (spi_data_out_r_39__N_1636[15]), 
            .\spi_data_out_r_39__N_1781[15] (spi_data_out_r_39__N_1781[15]), 
            .\spi_data_out_r_39__N_1636[14] (spi_data_out_r_39__N_1636[14]), 
            .\spi_data_out_r_39__N_1781[14] (spi_data_out_r_39__N_1781[14]), 
            .\spi_data_out_r_39__N_1636[13] (spi_data_out_r_39__N_1636[13]), 
            .\spi_data_out_r_39__N_1781[13] (spi_data_out_r_39__N_1781[13]), 
            .\spi_data_out_r_39__N_1636[12] (spi_data_out_r_39__N_1636[12]), 
            .\spi_data_out_r_39__N_1781[12] (spi_data_out_r_39__N_1781[12]), 
            .\spi_data_out_r_39__N_1636[11] (spi_data_out_r_39__N_1636[11]), 
            .\spi_data_out_r_39__N_1781[11] (spi_data_out_r_39__N_1781[11]), 
            .\spi_data_out_r_39__N_1636[10] (spi_data_out_r_39__N_1636[10]), 
            .\spi_data_out_r_39__N_1781[10] (spi_data_out_r_39__N_1781[10]), 
            .\spi_data_out_r_39__N_1636[9] (spi_data_out_r_39__N_1636[9]), 
            .\spi_data_out_r_39__N_1781[9] (spi_data_out_r_39__N_1781[9]), 
            .\spi_data_out_r_39__N_1636[8] (spi_data_out_r_39__N_1636[8]), 
            .\spi_data_out_r_39__N_1781[8] (spi_data_out_r_39__N_1781[8]), 
            .\spi_data_out_r_39__N_1636[7] (spi_data_out_r_39__N_1636[7]), 
            .\spi_data_out_r_39__N_1781[7] (spi_data_out_r_39__N_1781[7]), 
            .\spi_data_out_r_39__N_1636[6] (spi_data_out_r_39__N_1636[6]), 
            .\spi_data_out_r_39__N_1781[6] (spi_data_out_r_39__N_1781[6]), 
            .\spi_data_out_r_39__N_1636[5] (spi_data_out_r_39__N_1636[5]), 
            .\spi_data_out_r_39__N_1781[5] (spi_data_out_r_39__N_1781[5]), 
            .\spi_data_out_r_39__N_1636[4] (spi_data_out_r_39__N_1636[4]), 
            .\spi_data_out_r_39__N_1781[4] (spi_data_out_r_39__N_1781[4]), 
            .\spi_data_out_r_39__N_1636[3] (spi_data_out_r_39__N_1636[3]), 
            .\spi_data_out_r_39__N_1781[3] (spi_data_out_r_39__N_1781[3]), 
            .\spi_data_out_r_39__N_1636[2] (spi_data_out_r_39__N_1636[2]), 
            .\spi_data_out_r_39__N_1781[2] (spi_data_out_r_39__N_1781[2]), 
            .\spi_data_out_r_39__N_1636[1] (spi_data_out_r_39__N_1636[1]), 
            .\spi_data_out_r_39__N_1781[1] (spi_data_out_r_39__N_1781[1]), 
            .\spi_data_r[1] (spi_data_r[1]), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[3] (spi_data_r[3]), .\spi_data_r[4] (spi_data_r[4]), 
            .\spi_data_r[5] (spi_data_r[5]), .\spi_data_r[6] (spi_data_r[6]), 
            .\spi_data_r[7] (spi_data_r[7]), .\spi_data_r[8] (spi_data_r[8]), 
            .\spi_data_r[9] (spi_data_r[9]), .\spi_data_r[10] (spi_data_r[10]), 
            .\spi_data_r[11] (spi_data_r[11]), .\spi_data_r[12] (spi_data_r[12]), 
            .\spi_data_r[13] (spi_data_r[13]), .\spi_data_r[14] (spi_data_r[14]), 
            .\spi_data_r[15] (spi_data_r[15]), .\spi_data_r[16] (spi_data_r[16]), 
            .\spi_data_r[17] (spi_data_r[17]), .\spi_data_r[18] (spi_data_r[18]), 
            .\spi_data_r[19] (spi_data_r[19]), .\spi_data_r[20] (spi_data_r[20]), 
            .\spi_data_r[21] (spi_data_r[21]), .\spi_data_r[22] (spi_data_r[22]), 
            .\spi_data_r[23] (spi_data_r[23]), .\spi_data_r[24] (spi_data_r[24]), 
            .\spi_data_r[25] (spi_data_r[25]), .\spi_data_r[26] (spi_data_r[26]), 
            .\spi_data_r[27] (spi_data_r[27]), .\spi_data_r[28] (spi_data_r[28]), 
            .\spi_data_r[29] (spi_data_r[29]), .\spi_data_r[30] (spi_data_r[30]), 
            .\spi_data_r[31] (spi_data_r[31]), .\quad_homing[1] (quad_homing_adj_8343[1]), 
            .clk_enable_505(clk_enable_505), .n29120(n29120), .n13052(n13052), 
            .n26969(n26969), .pin_io_out_34(pin_io_out_34), .n27632(n27632)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(272[3] 293[2])
    \servo(DEV_ID=6,UART_ADDRESS_WIDTH=4)  \servo_ins_6..u_servo  (.mode(mode_adj_8127), 
            .clk(clk), .clk_enable_170(clk_enable_170), .n29239(n29239), 
            .\spi_data_r[0] (spi_data_r[0]), .n29191(n29191), .n29196(n29196), 
            .mode_adj_182(mode_adj_8124), .n14(n14), .C_5_c_c(C_5_c_c), 
            .n29267(n29267), .n8633(n8633)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(418[3] 453[2])
    \quad_decoder(DEV_ID=4)  \quad_ins_4..u_quad_decoder  (.quad_count({quad_count_adj_8403}), 
            .clk_1MHz(clk_1MHz), .\spi_data_out_r_39__N_1870[0] (spi_data_out_r_39__N_1870[0]), 
            .clk(clk), .\spi_data_out_r_39__N_2015[0] (spi_data_out_r_39__N_2015[0]), 
            .\quad_b[4] (quad_b[4]), .quad_buffer({quad_buffer_adj_8404}), 
            .\pin_intrpt[14] (pin_intrpt[14]), .n29239(n29239), .clk_enable_162(clk_enable_162), 
            .\spi_data_r[0] (spi_data_r[0]), .quad_homing({quad_homing_adj_8402}), 
            .clk_enable_77(clk_enable_77), .n29762(n29762), .\spi_data_r[1] (spi_data_r[1]), 
            .\spi_data_r[31] (spi_data_r[31]), .\spi_data_r[30] (spi_data_r[30]), 
            .\spi_data_r[29] (spi_data_r[29]), .\spi_data_r[28] (spi_data_r[28]), 
            .\spi_data_r[27] (spi_data_r[27]), .\spi_data_r[26] (spi_data_r[26]), 
            .\spi_data_r[25] (spi_data_r[25]), .\spi_data_r[24] (spi_data_r[24]), 
            .\spi_data_r[23] (spi_data_r[23]), .\spi_data_r[22] (spi_data_r[22]), 
            .\spi_data_r[21] (spi_data_r[21]), .\spi_data_r[20] (spi_data_r[20]), 
            .\spi_data_r[19] (spi_data_r[19]), .\spi_data_r[18] (spi_data_r[18]), 
            .\spi_data_r[17] (spi_data_r[17]), .\spi_data_r[16] (spi_data_r[16]), 
            .\spi_data_r[15] (spi_data_r[15]), .\spi_data_r[14] (spi_data_r[14]), 
            .\spi_data_r[13] (spi_data_r[13]), .\spi_data_r[12] (spi_data_r[12]), 
            .\spi_data_r[11] (spi_data_r[11]), .\spi_data_r[10] (spi_data_r[10]), 
            .\spi_data_r[9] (spi_data_r[9]), .\spi_data_r[8] (spi_data_r[8]), 
            .\spi_data_r[7] (spi_data_r[7]), .\spi_data_r[6] (spi_data_r[6]), 
            .\spi_data_r[5] (spi_data_r[5]), .\spi_data_r[4] (spi_data_r[4]), 
            .\spi_data_r[3] (spi_data_r[3]), .\spi_data_r[2] (spi_data_r[2]), 
            .quad_set_complete(quad_set_complete_adj_7757), .spi_data_out_r_39__N_1910(spi_data_out_r_39__N_1910), 
            .spi_data_out_r_39__N_2098(spi_data_out_r_39__N_2098), .\quad_a[4] (quad_a[4]), 
            .\spi_data_out_r_39__N_1870[31] (spi_data_out_r_39__N_1870[31]), 
            .\spi_data_out_r_39__N_2015[31] (spi_data_out_r_39__N_2015[31]), 
            .\spi_data_out_r_39__N_1870[30] (spi_data_out_r_39__N_1870[30]), 
            .\spi_data_out_r_39__N_2015[30] (spi_data_out_r_39__N_2015[30]), 
            .\spi_data_out_r_39__N_1870[29] (spi_data_out_r_39__N_1870[29]), 
            .\spi_data_out_r_39__N_2015[29] (spi_data_out_r_39__N_2015[29]), 
            .\spi_data_out_r_39__N_1870[28] (spi_data_out_r_39__N_1870[28]), 
            .\spi_data_out_r_39__N_2015[28] (spi_data_out_r_39__N_2015[28]), 
            .\spi_data_out_r_39__N_1870[27] (spi_data_out_r_39__N_1870[27]), 
            .\spi_data_out_r_39__N_2015[27] (spi_data_out_r_39__N_2015[27]), 
            .\spi_data_out_r_39__N_1870[26] (spi_data_out_r_39__N_1870[26]), 
            .\spi_data_out_r_39__N_2015[26] (spi_data_out_r_39__N_2015[26]), 
            .\spi_data_out_r_39__N_1870[25] (spi_data_out_r_39__N_1870[25]), 
            .\spi_data_out_r_39__N_2015[25] (spi_data_out_r_39__N_2015[25]), 
            .\spi_data_out_r_39__N_1870[24] (spi_data_out_r_39__N_1870[24]), 
            .\spi_data_out_r_39__N_2015[24] (spi_data_out_r_39__N_2015[24]), 
            .\spi_data_out_r_39__N_1870[23] (spi_data_out_r_39__N_1870[23]), 
            .\spi_data_out_r_39__N_2015[23] (spi_data_out_r_39__N_2015[23]), 
            .\spi_data_out_r_39__N_1870[22] (spi_data_out_r_39__N_1870[22]), 
            .\spi_data_out_r_39__N_2015[22] (spi_data_out_r_39__N_2015[22]), 
            .\spi_data_out_r_39__N_1870[21] (spi_data_out_r_39__N_1870[21]), 
            .\spi_data_out_r_39__N_2015[21] (spi_data_out_r_39__N_2015[21]), 
            .\spi_data_out_r_39__N_1870[20] (spi_data_out_r_39__N_1870[20]), 
            .\spi_data_out_r_39__N_2015[20] (spi_data_out_r_39__N_2015[20]), 
            .\spi_data_out_r_39__N_1870[19] (spi_data_out_r_39__N_1870[19]), 
            .\spi_data_out_r_39__N_2015[19] (spi_data_out_r_39__N_2015[19]), 
            .\spi_data_out_r_39__N_1870[18] (spi_data_out_r_39__N_1870[18]), 
            .\spi_data_out_r_39__N_2015[18] (spi_data_out_r_39__N_2015[18]), 
            .\spi_data_out_r_39__N_1870[17] (spi_data_out_r_39__N_1870[17]), 
            .\spi_data_out_r_39__N_2015[17] (spi_data_out_r_39__N_2015[17]), 
            .\spi_data_out_r_39__N_1870[16] (spi_data_out_r_39__N_1870[16]), 
            .\spi_data_out_r_39__N_2015[16] (spi_data_out_r_39__N_2015[16]), 
            .\spi_data_out_r_39__N_1870[15] (spi_data_out_r_39__N_1870[15]), 
            .\spi_data_out_r_39__N_2015[15] (spi_data_out_r_39__N_2015[15]), 
            .\spi_data_out_r_39__N_1870[14] (spi_data_out_r_39__N_1870[14]), 
            .\spi_data_out_r_39__N_2015[14] (spi_data_out_r_39__N_2015[14]), 
            .\spi_data_out_r_39__N_1870[13] (spi_data_out_r_39__N_1870[13]), 
            .\spi_data_out_r_39__N_2015[13] (spi_data_out_r_39__N_2015[13]), 
            .\spi_data_out_r_39__N_1870[12] (spi_data_out_r_39__N_1870[12]), 
            .\spi_data_out_r_39__N_2015[12] (spi_data_out_r_39__N_2015[12]), 
            .\spi_data_out_r_39__N_1870[11] (spi_data_out_r_39__N_1870[11]), 
            .\spi_data_out_r_39__N_2015[11] (spi_data_out_r_39__N_2015[11]), 
            .\spi_data_out_r_39__N_1870[10] (spi_data_out_r_39__N_1870[10]), 
            .\spi_data_out_r_39__N_2015[10] (spi_data_out_r_39__N_2015[10]), 
            .\spi_data_out_r_39__N_1870[9] (spi_data_out_r_39__N_1870[9]), 
            .\spi_data_out_r_39__N_2015[9] (spi_data_out_r_39__N_2015[9]), 
            .\spi_data_out_r_39__N_1870[8] (spi_data_out_r_39__N_1870[8]), 
            .\spi_data_out_r_39__N_2015[8] (spi_data_out_r_39__N_2015[8]), 
            .\spi_data_out_r_39__N_1870[7] (spi_data_out_r_39__N_1870[7]), 
            .\spi_data_out_r_39__N_2015[7] (spi_data_out_r_39__N_2015[7]), 
            .\spi_data_out_r_39__N_1870[6] (spi_data_out_r_39__N_1870[6]), 
            .\spi_data_out_r_39__N_2015[6] (spi_data_out_r_39__N_2015[6]), 
            .\spi_data_out_r_39__N_1870[5] (spi_data_out_r_39__N_1870[5]), 
            .\spi_data_out_r_39__N_2015[5] (spi_data_out_r_39__N_2015[5]), 
            .\spi_data_out_r_39__N_1870[4] (spi_data_out_r_39__N_1870[4]), 
            .\spi_data_out_r_39__N_2015[4] (spi_data_out_r_39__N_2015[4]), 
            .\spi_data_out_r_39__N_1870[3] (spi_data_out_r_39__N_1870[3]), 
            .\spi_data_out_r_39__N_2015[3] (spi_data_out_r_39__N_2015[3]), 
            .\spi_data_out_r_39__N_1870[2] (spi_data_out_r_39__N_1870[2]), 
            .\spi_data_out_r_39__N_2015[2] (spi_data_out_r_39__N_2015[2]), 
            .\spi_data_out_r_39__N_1870[1] (spi_data_out_r_39__N_1870[1]), 
            .\spi_data_out_r_39__N_2015[1] (spi_data_out_r_39__N_2015[1]), 
            .resetn_c(resetn_c), .GND_net(GND_net), .clk_enable_518(clk_enable_518), 
            .n29080(n29080), .n26938(n26938)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(272[3] 293[2])
    \quad_decoder(DEV_ID=1)  \quad_ins_1..u_quad_decoder  (.clk(clk), .clk_enable_286(clk_enable_286), 
            .n29239(n29239), .n29762(n29762), .quad_count({quad_count_adj_8226}), 
            .clk_1MHz(clk_1MHz), .\spi_data_out_r_39__N_1168[0] (spi_data_out_r_39__N_1168[0]), 
            .\spi_data_out_r_39__N_1313[0] (spi_data_out_r_39__N_1313[0]), 
            .\quad_b[1] (quad_b[1]), .quad_buffer({quad_buffer_adj_8227}), 
            .\pin_intrpt[5] (pin_intrpt[5]), .clk_enable_467(clk_enable_467), 
            .\spi_data_r[0] (spi_data_r[0]), .quad_set_complete(quad_set_complete_adj_7619), 
            .spi_data_out_r_39__N_1208(spi_data_out_r_39__N_1208), .spi_data_out_r_39__N_1396(spi_data_out_r_39__N_1396), 
            .resetn_c(resetn_c), .GND_net(GND_net), .\quad_a[1] (quad_a[1]), 
            .\spi_data_out_r_39__N_1168[31] (spi_data_out_r_39__N_1168[31]), 
            .\spi_data_out_r_39__N_1313[31] (spi_data_out_r_39__N_1313[31]), 
            .\spi_data_out_r_39__N_1168[30] (spi_data_out_r_39__N_1168[30]), 
            .\spi_data_out_r_39__N_1313[30] (spi_data_out_r_39__N_1313[30]), 
            .\spi_data_out_r_39__N_1168[29] (spi_data_out_r_39__N_1168[29]), 
            .\spi_data_out_r_39__N_1313[29] (spi_data_out_r_39__N_1313[29]), 
            .\spi_data_out_r_39__N_1168[28] (spi_data_out_r_39__N_1168[28]), 
            .\spi_data_out_r_39__N_1313[28] (spi_data_out_r_39__N_1313[28]), 
            .\spi_data_out_r_39__N_1168[27] (spi_data_out_r_39__N_1168[27]), 
            .\spi_data_out_r_39__N_1313[27] (spi_data_out_r_39__N_1313[27]), 
            .\spi_data_out_r_39__N_1168[26] (spi_data_out_r_39__N_1168[26]), 
            .\spi_data_out_r_39__N_1313[26] (spi_data_out_r_39__N_1313[26]), 
            .\spi_data_out_r_39__N_1168[25] (spi_data_out_r_39__N_1168[25]), 
            .\spi_data_out_r_39__N_1313[25] (spi_data_out_r_39__N_1313[25]), 
            .\spi_data_out_r_39__N_1168[24] (spi_data_out_r_39__N_1168[24]), 
            .\spi_data_out_r_39__N_1313[24] (spi_data_out_r_39__N_1313[24]), 
            .\spi_data_out_r_39__N_1168[23] (spi_data_out_r_39__N_1168[23]), 
            .\spi_data_out_r_39__N_1313[23] (spi_data_out_r_39__N_1313[23]), 
            .\spi_data_out_r_39__N_1168[22] (spi_data_out_r_39__N_1168[22]), 
            .\spi_data_out_r_39__N_1313[22] (spi_data_out_r_39__N_1313[22]), 
            .\spi_data_out_r_39__N_1168[21] (spi_data_out_r_39__N_1168[21]), 
            .\spi_data_out_r_39__N_1313[21] (spi_data_out_r_39__N_1313[21]), 
            .\spi_data_out_r_39__N_1168[20] (spi_data_out_r_39__N_1168[20]), 
            .\spi_data_out_r_39__N_1313[20] (spi_data_out_r_39__N_1313[20]), 
            .\spi_data_out_r_39__N_1168[19] (spi_data_out_r_39__N_1168[19]), 
            .\spi_data_out_r_39__N_1313[19] (spi_data_out_r_39__N_1313[19]), 
            .\spi_data_out_r_39__N_1168[18] (spi_data_out_r_39__N_1168[18]), 
            .\spi_data_out_r_39__N_1313[18] (spi_data_out_r_39__N_1313[18]), 
            .\spi_data_out_r_39__N_1168[17] (spi_data_out_r_39__N_1168[17]), 
            .\spi_data_out_r_39__N_1313[17] (spi_data_out_r_39__N_1313[17]), 
            .\spi_data_out_r_39__N_1168[16] (spi_data_out_r_39__N_1168[16]), 
            .\spi_data_out_r_39__N_1313[16] (spi_data_out_r_39__N_1313[16]), 
            .\spi_data_out_r_39__N_1168[15] (spi_data_out_r_39__N_1168[15]), 
            .\spi_data_out_r_39__N_1313[15] (spi_data_out_r_39__N_1313[15]), 
            .\spi_data_out_r_39__N_1168[14] (spi_data_out_r_39__N_1168[14]), 
            .\spi_data_out_r_39__N_1313[14] (spi_data_out_r_39__N_1313[14]), 
            .\spi_data_out_r_39__N_1168[13] (spi_data_out_r_39__N_1168[13]), 
            .\spi_data_out_r_39__N_1313[13] (spi_data_out_r_39__N_1313[13]), 
            .\spi_data_out_r_39__N_1168[12] (spi_data_out_r_39__N_1168[12]), 
            .\spi_data_out_r_39__N_1313[12] (spi_data_out_r_39__N_1313[12]), 
            .\spi_data_out_r_39__N_1168[11] (spi_data_out_r_39__N_1168[11]), 
            .\spi_data_out_r_39__N_1313[11] (spi_data_out_r_39__N_1313[11]), 
            .\spi_data_out_r_39__N_1168[10] (spi_data_out_r_39__N_1168[10]), 
            .\spi_data_out_r_39__N_1313[10] (spi_data_out_r_39__N_1313[10]), 
            .\spi_data_out_r_39__N_1168[9] (spi_data_out_r_39__N_1168[9]), 
            .\spi_data_out_r_39__N_1313[9] (spi_data_out_r_39__N_1313[9]), 
            .\spi_data_out_r_39__N_1168[8] (spi_data_out_r_39__N_1168[8]), 
            .\spi_data_out_r_39__N_1313[8] (spi_data_out_r_39__N_1313[8]), 
            .\spi_data_out_r_39__N_1168[7] (spi_data_out_r_39__N_1168[7]), 
            .\spi_data_out_r_39__N_1313[7] (spi_data_out_r_39__N_1313[7]), 
            .\spi_data_out_r_39__N_1168[6] (spi_data_out_r_39__N_1168[6]), 
            .\spi_data_out_r_39__N_1313[6] (spi_data_out_r_39__N_1313[6]), 
            .\spi_data_out_r_39__N_1168[5] (spi_data_out_r_39__N_1168[5]), 
            .\spi_data_out_r_39__N_1313[5] (spi_data_out_r_39__N_1313[5]), 
            .\spi_data_out_r_39__N_1168[4] (spi_data_out_r_39__N_1168[4]), 
            .\spi_data_out_r_39__N_1313[4] (spi_data_out_r_39__N_1313[4]), 
            .\spi_data_out_r_39__N_1168[3] (spi_data_out_r_39__N_1168[3]), 
            .\spi_data_out_r_39__N_1313[3] (spi_data_out_r_39__N_1313[3]), 
            .\spi_data_out_r_39__N_1168[2] (spi_data_out_r_39__N_1168[2]), 
            .\spi_data_out_r_39__N_1313[2] (spi_data_out_r_39__N_1313[2]), 
            .\spi_data_out_r_39__N_1168[1] (spi_data_out_r_39__N_1168[1]), 
            .\spi_data_out_r_39__N_1313[1] (spi_data_out_r_39__N_1313[1]), 
            .\quad_homing[1] (quad_homing_adj_8225[1]), .\spi_data_r[1] (spi_data_r[1]), 
            .\spi_data_r[2] (spi_data_r[2]), .\spi_data_r[3] (spi_data_r[3]), 
            .\spi_data_r[4] (spi_data_r[4]), .\spi_data_r[5] (spi_data_r[5]), 
            .\spi_data_r[6] (spi_data_r[6]), .\spi_data_r[7] (spi_data_r[7]), 
            .\spi_data_r[8] (spi_data_r[8]), .\spi_data_r[9] (spi_data_r[9]), 
            .\spi_data_r[10] (spi_data_r[10]), .\spi_data_r[11] (spi_data_r[11]), 
            .\spi_data_r[12] (spi_data_r[12]), .\spi_data_r[13] (spi_data_r[13]), 
            .\spi_data_r[14] (spi_data_r[14]), .\spi_data_r[15] (spi_data_r[15]), 
            .\spi_data_r[16] (spi_data_r[16]), .\spi_data_r[17] (spi_data_r[17]), 
            .\spi_data_r[18] (spi_data_r[18]), .\spi_data_r[19] (spi_data_r[19]), 
            .\spi_data_r[20] (spi_data_r[20]), .\spi_data_r[21] (spi_data_r[21]), 
            .\spi_data_r[22] (spi_data_r[22]), .\spi_data_r[23] (spi_data_r[23]), 
            .\spi_data_r[24] (spi_data_r[24]), .\spi_data_r[25] (spi_data_r[25]), 
            .\spi_data_r[26] (spi_data_r[26]), .\spi_data_r[27] (spi_data_r[27]), 
            .\spi_data_r[28] (spi_data_r[28]), .\spi_data_r[29] (spi_data_r[29]), 
            .\spi_data_r[30] (spi_data_r[30]), .\spi_data_r[31] (spi_data_r[31]), 
            .clk_enable_502(clk_enable_502), .n29084(n29084), .n12716(n12716), 
            .n26963(n26963), .pin_io_out_14(pin_io_out_14), .n27636(n27636)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(272[3] 293[2])
    \stepper(DEV_ID=6,UART_ADDRESS_WIDTH=4)  \stepper_ins_6..u_stepper  (.\spi_data_out_r[26] (spi_data_out_r[26]), 
            .\spi_data_out_r_39__N_1168[26] (spi_data_out_r_39__N_1168[26]), 
            .spi_data_out_r_39__N_1208(spi_data_out_r_39__N_1208), .mode_adj_181({n29786}), 
            .clk(clk), .clk_enable_288(clk_enable_288), .n29239(n29239), 
            .n29762(n29762), .\spi_data_out_r_39__N_1636[15] (spi_data_out_r_39__N_1636[15]), 
            .spi_data_out_r_39__N_1676(spi_data_out_r_39__N_1676), .\spi_data_out_r_39__N_4835[26] (spi_data_out_r_39__N_4835[26]), 
            .spi_data_out_r_39__N_4875(spi_data_out_r_39__N_4875), .\spi_data_out_r_39__N_5513[26] (spi_data_out_r_39__N_5513[26]), 
            .spi_data_out_r_39__N_5553(spi_data_out_r_39__N_5553), .\spi_data_out_r_39__N_4496[26] (spi_data_out_r_39__N_4496[26]), 
            .spi_data_out_r_39__N_4536(spi_data_out_r_39__N_4536), .\spi_data_out_r_39__N_3818[26] (spi_data_out_r_39__N_3818[26]), 
            .spi_data_out_r_39__N_3858(spi_data_out_r_39__N_3858), .\spi_data_out_r_39__N_2104[26] (spi_data_out_r_39__N_2104[26]), 
            .\spi_data_out_r_39__N_1870[26] (spi_data_out_r_39__N_1870[26]), 
            .spi_data_out_r_39__N_2144(spi_data_out_r_39__N_2144), .spi_data_out_r_39__N_1910(spi_data_out_r_39__N_1910), 
            .\spi_data_out_r_39__N_1402[26] (spi_data_out_r_39__N_1402[26]), 
            .spi_data_out_r_39__N_1442(spi_data_out_r_39__N_1442), .\spi_data_out_r_39__N_2338[26] (spi_data_out_r_39__N_2338[26]), 
            .\spi_data_out_r_39__N_5174[26] (spi_data_out_r_39__N_5174[26]), 
            .spi_data_out_r_39__N_2378(spi_data_out_r_39__N_2378), .spi_data_out_r_39__N_5214(spi_data_out_r_39__N_5214), 
            .\spi_data_out_r_39__N_1636[26] (spi_data_out_r_39__N_1636[26]), 
            .\spi_data_out_r_39__N_934[26] (spi_data_out_r_39__N_934[26]), 
            .spi_data_out_r_39__N_974(spi_data_out_r_39__N_974), .spi_data_out_r_39__N_5892(spi_data_out_r_39__N_5892), 
            .\spi_data_out_r_39__N_4157[26] (spi_data_out_r_39__N_4157[26]), 
            .spi_data_out_r_39__N_4197(spi_data_out_r_39__N_4197), .pin_io_out_68(pin_io_out_68), 
            .\quad_a[6] (quad_a[6]), .n28811(n28811), .\spi_data_out_r[27] (spi_data_out_r[27]), 
            .pin_io_out_69(pin_io_out_69), .\quad_b[6] (quad_b[6]), .\spi_data_out_r_39__N_1168[27] (spi_data_out_r_39__N_1168[27]), 
            .\spi_data_out_r_39__N_4835[27] (spi_data_out_r_39__N_4835[27]), 
            .\spi_data_out_r_39__N_5513[27] (spi_data_out_r_39__N_5513[27]), 
            .\spi_data_out_r_39__N_4835[21] (spi_data_out_r_39__N_4835[21]), 
            .\spi_data_out_r_39__N_4496[27] (spi_data_out_r_39__N_4496[27]), 
            .\spi_data_out_r_39__N_3818[27] (spi_data_out_r_39__N_3818[27]), 
            .\spi_data_out_r_39__N_2104[27] (spi_data_out_r_39__N_2104[27]), 
            .\spi_data_out_r_39__N_1870[27] (spi_data_out_r_39__N_1870[27]), 
            .\spi_data_out_r_39__N_1402[27] (spi_data_out_r_39__N_1402[27]), 
            .\spi_data_out_r_39__N_2338[27] (spi_data_out_r_39__N_2338[27]), 
            .\spi_data_out_r_39__N_5174[27] (spi_data_out_r_39__N_5174[27]), 
            .\spi_data_out_r_39__N_1636[27] (spi_data_out_r_39__N_1636[27]), 
            .\spi_data_out_r_39__N_934[27] (spi_data_out_r_39__N_934[27]), 
            .\spi_data_out_r_39__N_4157[27] (spi_data_out_r_39__N_4157[27]), 
            .\spi_data_out_r[28] (spi_data_out_r[28]), .\spi_data_out_r_39__N_1168[28] (spi_data_out_r_39__N_1168[28]), 
            .\SLO_buf[0] (SLO_buf_adj_8951[0]), .\spi_data_out_r_39__N_5852[0] (spi_data_out_r_39__N_5852[0]), 
            .\spi_data_out_r_39__N_6114[0] (spi_data_out_r_39__N_6114[0]), 
            .\spi_data_out_r_39__N_4835[28] (spi_data_out_r_39__N_4835[28]), 
            .clk_1MHz(clk_1MHz), .clk_1MHz_enable_367(clk_1MHz_enable_367), 
            .\spi_data_out_r_39__N_5513[28] (spi_data_out_r_39__N_5513[28]), 
            .\spi_data_out_r_39__N_934[15] (spi_data_out_r_39__N_934[15]), 
            .\spi_data_out_r_39__N_4157[15] (spi_data_out_r_39__N_4157[15]), 
            .\spi_data_out_r_39__N_4496[28] (spi_data_out_r_39__N_4496[28]), 
            .\spi_data_out_r_39__N_3818[28] (spi_data_out_r_39__N_3818[28]), 
            .\spi_data_out_r_39__N_2104[28] (spi_data_out_r_39__N_2104[28]), 
            .\spi_data_out_r_39__N_1870[28] (spi_data_out_r_39__N_1870[28]), 
            .\spi_data_out_r_39__N_1402[28] (spi_data_out_r_39__N_1402[28]), 
            .\spi_data_out_r_39__N_2338[28] (spi_data_out_r_39__N_2338[28]), 
            .\spi_data_out_r_39__N_5174[28] (spi_data_out_r_39__N_5174[28]), 
            .\spi_data_out_r_39__N_1636[21] (spi_data_out_r_39__N_1636[21]), 
            .\spi_data_out_r_39__N_934[21] (spi_data_out_r_39__N_934[21]), 
            .\spi_data_out_r_39__N_4157[21] (spi_data_out_r_39__N_4157[21]), 
            .\spi_data_out_r_39__N_1636[28] (spi_data_out_r_39__N_1636[28]), 
            .\spi_data_out_r[22] (spi_data_out_r[22]), .\spi_data_out_r_39__N_1168[22] (spi_data_out_r_39__N_1168[22]), 
            .\spi_data_out_r_39__N_4835[22] (spi_data_out_r_39__N_4835[22]), 
            .\spi_data_out_r_39__N_5513[22] (spi_data_out_r_39__N_5513[22]), 
            .\spi_data_out_r_39__N_934[28] (spi_data_out_r_39__N_934[28]), 
            .\spi_data_out_r_39__N_4157[28] (spi_data_out_r_39__N_4157[28]), 
            .\spi_data_out_r[29] (spi_data_out_r[29]), .\spi_data_out_r_39__N_4496[22] (spi_data_out_r_39__N_4496[22]), 
            .\spi_data_out_r_39__N_1168[29] (spi_data_out_r_39__N_1168[29]), 
            .\spi_data_out_r_39__N_4835[29] (spi_data_out_r_39__N_4835[29]), 
            .\spi_data_out_r_39__N_5513[29] (spi_data_out_r_39__N_5513[29]), 
            .\spi_data_out_r_39__N_4496[29] (spi_data_out_r_39__N_4496[29]), 
            .\spi_data_out_r_39__N_3818[29] (spi_data_out_r_39__N_3818[29]), 
            .\spi_data_out_r_39__N_3818[22] (spi_data_out_r_39__N_3818[22]), 
            .\spi_data_out_r_39__N_2104[29] (spi_data_out_r_39__N_2104[29]), 
            .\spi_data_out_r_39__N_1870[29] (spi_data_out_r_39__N_1870[29]), 
            .\spi_data_out_r_39__N_2104[22] (spi_data_out_r_39__N_2104[22]), 
            .\spi_data_out_r_39__N_1870[22] (spi_data_out_r_39__N_1870[22]), 
            .\spi_data_out_r_39__N_1402[22] (spi_data_out_r_39__N_1402[22]), 
            .\spi_data_out_r_39__N_1402[29] (spi_data_out_r_39__N_1402[29]), 
            .\spi_data_out_r_39__N_2338[29] (spi_data_out_r_39__N_2338[29]), 
            .\spi_data_out_r_39__N_5174[29] (spi_data_out_r_39__N_5174[29]), 
            .\spi_data_out_r_39__N_1636[29] (spi_data_out_r_39__N_1636[29]), 
            .\spi_data_out_r_39__N_2338[22] (spi_data_out_r_39__N_2338[22]), 
            .\spi_data_out_r_39__N_5174[22] (spi_data_out_r_39__N_5174[22]), 
            .\spi_data_out_r_39__N_934[29] (spi_data_out_r_39__N_934[29]), 
            .n29087(n29087), .\spi_data_out_r_39__N_4157[29] (spi_data_out_r_39__N_4157[29]), 
            .\spi_data_out_r_39__N_1636[22] (spi_data_out_r_39__N_1636[22]), 
            .\spi_data_out_r[30] (spi_data_out_r[30]), .\spi_data_out_r_39__N_1168[30] (spi_data_out_r_39__N_1168[30]), 
            .\spi_data_out_r_39__N_934[22] (spi_data_out_r_39__N_934[22]), 
            .\spi_data_out_r_39__N_4835[30] (spi_data_out_r_39__N_4835[30]), 
            .\spi_data_out_r_39__N_5513[30] (spi_data_out_r_39__N_5513[30]), 
            .\spi_data_out_r_39__N_4157[22] (spi_data_out_r_39__N_4157[22]), 
            .\spi_data_out_r_39__N_4496[30] (spi_data_out_r_39__N_4496[30]), 
            .\spi_data_out_r[23] (spi_data_out_r[23]), .\spi_data_out_r_39__N_3818[30] (spi_data_out_r_39__N_3818[30]), 
            .digital_output_r(digital_output_r_adj_8090), .clk_enable_198(clk_enable_198), 
            .\spi_data_r[0] (spi_data_r[0]), .\spi_data_out_r_39__N_1168[23] (spi_data_out_r_39__N_1168[23]), 
            .\spi_data_out_r_39__N_2104[30] (spi_data_out_r_39__N_2104[30]), 
            .\spi_data_out_r_39__N_1870[30] (spi_data_out_r_39__N_1870[30]), 
            .\spi_data_out_r_39__N_1402[30] (spi_data_out_r_39__N_1402[30]), 
            .\spi_data_out_r_39__N_2338[30] (spi_data_out_r_39__N_2338[30]), 
            .\spi_data_out_r_39__N_5174[30] (spi_data_out_r_39__N_5174[30]), 
            .\spi_data_out_r_39__N_1636[30] (spi_data_out_r_39__N_1636[30]), 
            .\spi_data_out_r_39__N_934[30] (spi_data_out_r_39__N_934[30]), 
            .\spi_data_out_r_39__N_4157[30] (spi_data_out_r_39__N_4157[30]), 
            .\spi_data_out_r[31] (spi_data_out_r[31]), .\spi_data_out_r_39__N_4835[23] (spi_data_out_r_39__N_4835[23]), 
            .\spi_data_out_r_39__N_1168[31] (spi_data_out_r_39__N_1168[31]), 
            .\spi_data_out_r_39__N_5513[23] (spi_data_out_r_39__N_5513[23]), 
            .\spi_data_out_r[16] (spi_data_out_r[16]), .\spi_data_out_r_39__N_1168[16] (spi_data_out_r_39__N_1168[16]), 
            .\spi_data_out_r_39__N_4496[23] (spi_data_out_r_39__N_4496[23]), 
            .\spi_data_out_r_39__N_4835[31] (spi_data_out_r_39__N_4835[31]), 
            .\spi_data_out_r_39__N_3818[23] (spi_data_out_r_39__N_3818[23]), 
            .\spi_data_out_r_39__N_5513[31] (spi_data_out_r_39__N_5513[31]), 
            .\spi_data_out_r_39__N_4496[31] (spi_data_out_r_39__N_4496[31]), 
            .n19401(n19401), .resetn_c(resetn_c), .\spi_data_out_r_39__N_3818[31] (spi_data_out_r_39__N_3818[31]), 
            .\spi_data_out_r_39__N_2104[31] (spi_data_out_r_39__N_2104[31]), 
            .\spi_data_out_r_39__N_1870[31] (spi_data_out_r_39__N_1870[31]), 
            .\spi_data_out_r_39__N_1402[31] (spi_data_out_r_39__N_1402[31]), 
            .\spi_data_out_r_39__N_2338[31] (spi_data_out_r_39__N_2338[31]), 
            .\spi_data_out_r_39__N_5174[31] (spi_data_out_r_39__N_5174[31]), 
            .\spi_data_out_r_39__N_1636[31] (spi_data_out_r_39__N_1636[31]), 
            .\spi_data_out_r_39__N_934[31] (spi_data_out_r_39__N_934[31]), 
            .\spi_data_out_r_39__N_4157[31] (spi_data_out_r_39__N_4157[31]), 
            .\spi_data_out_r_39__N_4835[32] (spi_data_out_r_39__N_4835[32]), 
            .\spi_data_out_r[32] (spi_data_out_r[32]), .\spi_data_out_r_39__N_3818[32] (spi_data_out_r_39__N_3818[32]), 
            .\spi_data_out_r_39__N_5174[32] (spi_data_out_r_39__N_5174[32]), 
            .\spi_data_out_r_39__N_4496[32] (spi_data_out_r_39__N_4496[32]), 
            .\spi_data_out_r_39__N_4157[32] (spi_data_out_r_39__N_4157[32]), 
            .\spi_data_out_r_39__N_5513[32] (spi_data_out_r_39__N_5513[32]), 
            .\spi_data_out_r_39__N_4835[33] (spi_data_out_r_39__N_4835[33]), 
            .\spi_data_out_r[33] (spi_data_out_r[33]), .\spi_data_out_r_39__N_3818[33] (spi_data_out_r_39__N_3818[33]), 
            .\spi_data_out_r_39__N_5174[33] (spi_data_out_r_39__N_5174[33]), 
            .\spi_data_out_r_39__N_4496[33] (spi_data_out_r_39__N_4496[33]), 
            .\spi_data_out_r_39__N_4157[33] (spi_data_out_r_39__N_4157[33]), 
            .\spi_data_out_r_39__N_5513[33] (spi_data_out_r_39__N_5513[33]), 
            .\spi_data_out_r_39__N_4835[34] (spi_data_out_r_39__N_4835[34]), 
            .\spi_data_out_r[34] (spi_data_out_r[34]), .\spi_data_out_r_39__N_3818[34] (spi_data_out_r_39__N_3818[34]), 
            .\spi_data_out_r_39__N_5174[34] (spi_data_out_r_39__N_5174[34]), 
            .\spi_data_out_r_39__N_4496[34] (spi_data_out_r_39__N_4496[34]), 
            .\spi_data_out_r_39__N_4157[34] (spi_data_out_r_39__N_4157[34]), 
            .\spi_data_out_r_39__N_2104[23] (spi_data_out_r_39__N_2104[23]), 
            .\spi_data_out_r_39__N_1870[23] (spi_data_out_r_39__N_1870[23]), 
            .\spi_data_out_r_39__N_5513[34] (spi_data_out_r_39__N_5513[34]), 
            .\spi_data_out_r_39__N_4835[35] (spi_data_out_r_39__N_4835[35]), 
            .\spi_data_out_r[35] (spi_data_out_r[35]), .\spi_data_out_r_39__N_3818[35] (spi_data_out_r_39__N_3818[35]), 
            .\spi_data_out_r_39__N_5174[35] (spi_data_out_r_39__N_5174[35]), 
            .\spi_data_out_r_39__N_4496[35] (spi_data_out_r_39__N_4496[35]), 
            .\spi_data_out_r_39__N_4157[35] (spi_data_out_r_39__N_4157[35]), 
            .\spi_data_out_r_39__N_5513[35] (spi_data_out_r_39__N_5513[35]), 
            .\spi_data_out_r_39__N_4835[36] (spi_data_out_r_39__N_4835[36]), 
            .\spi_data_out_r[36] (spi_data_out_r[36]), .\spi_data_out_r_39__N_3818[36] (spi_data_out_r_39__N_3818[36]), 
            .\spi_data_out_r_39__N_5174[36] (spi_data_out_r_39__N_5174[36]), 
            .\spi_data_out_r_39__N_4496[36] (spi_data_out_r_39__N_4496[36]), 
            .\spi_data_out_r_39__N_4157[36] (spi_data_out_r_39__N_4157[36]), 
            .\spi_data_out_r_39__N_5513[36] (spi_data_out_r_39__N_5513[36]), 
            .\spi_data_out_r_39__N_4835[37] (spi_data_out_r_39__N_4835[37]), 
            .\spi_data_out_r[37] (spi_data_out_r[37]), .\spi_data_out_r_39__N_1402[23] (spi_data_out_r_39__N_1402[23]), 
            .\spi_data_out_r_39__N_3818[37] (spi_data_out_r_39__N_3818[37]), 
            .\spi_data_out_r_39__N_5174[37] (spi_data_out_r_39__N_5174[37]), 
            .\spi_data_out_r_39__N_4496[37] (spi_data_out_r_39__N_4496[37]), 
            .\spi_data_out_r_39__N_4157[37] (spi_data_out_r_39__N_4157[37]), 
            .\spi_data_out_r_39__N_2338[23] (spi_data_out_r_39__N_2338[23]), 
            .\spi_data_out_r_39__N_5174[23] (spi_data_out_r_39__N_5174[23]), 
            .\spi_data_out_r_39__N_5513[37] (spi_data_out_r_39__N_5513[37]), 
            .\spi_data_out_r_39__N_4835[38] (spi_data_out_r_39__N_4835[38]), 
            .\spi_data_out_r[38] (spi_data_out_r[38]), .\spi_data_out_r_39__N_3818[38] (spi_data_out_r_39__N_3818[38]), 
            .\spi_data_out_r_39__N_1636[23] (spi_data_out_r_39__N_1636[23]), 
            .\spi_data_out_r_39__N_5174[38] (spi_data_out_r_39__N_5174[38]), 
            .\spi_data_out_r_39__N_4496[38] (spi_data_out_r_39__N_4496[38]), 
            .\spi_data_out_r_39__N_4157[38] (spi_data_out_r_39__N_4157[38]), 
            .\spi_data_out_r_39__N_934[23] (spi_data_out_r_39__N_934[23]), 
            .\spi_data_out_r_39__N_4157[23] (spi_data_out_r_39__N_4157[23]), 
            .\spi_data_out_r_39__N_5513[38] (spi_data_out_r_39__N_5513[38]), 
            .\spi_data_out_r_39__N_4835[39] (spi_data_out_r_39__N_4835[39]), 
            .\spi_data_out_r[39] (spi_data_out_r[39]), .\spi_data_out_r_39__N_3818[39] (spi_data_out_r_39__N_3818[39]), 
            .\spi_data_out_r_39__N_5174[39] (spi_data_out_r_39__N_5174[39]), 
            .\spi_data_out_r_39__N_4496[39] (spi_data_out_r_39__N_4496[39]), 
            .\spi_data_out_r_39__N_4157[39] (spi_data_out_r_39__N_4157[39]), 
            .\spi_data_out_r_39__N_5513[39] (spi_data_out_r_39__N_5513[39]), 
            .\spi_data_out_r[24] (spi_data_out_r[24]), .\spi_data_out_r_39__N_1168[24] (spi_data_out_r_39__N_1168[24]), 
            .\spi_data_out_r_39__N_4835[24] (spi_data_out_r_39__N_4835[24]), 
            .\spi_data_out_r_39__N_5513[24] (spi_data_out_r_39__N_5513[24]), 
            .\spi_data_out_r_39__N_4496[24] (spi_data_out_r_39__N_4496[24]), 
            .n29267(n29267), .mode(mode_adj_8150), .n29191(n29191), .n29153(n29153), 
            .\spi_data_out_r_39__N_3818[24] (spi_data_out_r_39__N_3818[24]), 
            .n29195(n29195), .\spi_data_out_r_39__N_2104[24] (spi_data_out_r_39__N_2104[24]), 
            .\spi_data_out_r_39__N_1870[24] (spi_data_out_r_39__N_1870[24]), 
            .n29293(n29293), .\cs_decoded[12] (cs_decoded[12]), .n8652(n8652), 
            .n1(n1_adj_8154), .n8651(n8651), .n1_adj_171(n1), .\spi_data_out_r_39__N_5513[21] (spi_data_out_r_39__N_5513[21]), 
            .\spi_data_out_r_39__N_1402[24] (spi_data_out_r_39__N_1402[24]), 
            .\spi_data_out_r_39__N_2338[24] (spi_data_out_r_39__N_2338[24]), 
            .\spi_data_out_r_39__N_5174[24] (spi_data_out_r_39__N_5174[24]), 
            .\spi_data_out_r_39__N_1636[24] (spi_data_out_r_39__N_1636[24]), 
            .\spi_data_out_r_39__N_934[24] (spi_data_out_r_39__N_934[24]), 
            .\spi_data_out_r_39__N_4157[24] (spi_data_out_r_39__N_4157[24]), 
            .\spi_data_out_r[25] (spi_data_out_r[25]), .\spi_data_out_r_39__N_1168[25] (spi_data_out_r_39__N_1168[25]), 
            .\spi_data_out_r_39__N_4835[25] (spi_data_out_r_39__N_4835[25]), 
            .\spi_data_out_r_39__N_5513[25] (spi_data_out_r_39__N_5513[25]), 
            .\spi_data_out_r_39__N_4496[25] (spi_data_out_r_39__N_4496[25]), 
            .\spi_data_out_r_39__N_3818[25] (spi_data_out_r_39__N_3818[25]), 
            .\spi_data_out_r_39__N_2104[25] (spi_data_out_r_39__N_2104[25]), 
            .\spi_data_out_r_39__N_1870[25] (spi_data_out_r_39__N_1870[25]), 
            .\spi_data_out_r_39__N_1402[25] (spi_data_out_r_39__N_1402[25]), 
            .\spi_data_out_r_39__N_2338[25] (spi_data_out_r_39__N_2338[25]), 
            .\spi_data_out_r_39__N_5174[25] (spi_data_out_r_39__N_5174[25]), 
            .GND_net(GND_net), .\spi_data_out_r_39__N_1636[25] (spi_data_out_r_39__N_1636[25]), 
            .\spi_data_out_r_39__N_934[25] (spi_data_out_r_39__N_934[25]), 
            .\spi_data_out_r_39__N_4157[25] (spi_data_out_r_39__N_4157[25]), 
            .\spi_data_r[2] (spi_data_r[2]), .\spi_data_r[1] (spi_data_r[1]), 
            .\spi_data_out_r_39__N_4835[16] (spi_data_out_r_39__N_4835[16]), 
            .\spi_data_out_r_39__N_2856[2] (spi_data_out_r_39__N_2856[2]), 
            .clear_intrpt(clear_intrpt_adj_7960), .n13(n13), .\spi_data_out_r_39__N_1402[2] (spi_data_out_r_39__N_1402[2]), 
            .n4(n4), .\SLO_buf[1] (SLO_buf_adj_8951[1]), .\SLO_buf[2] (SLO_buf_adj_8951[2]), 
            .\SLO_buf[3] (SLO_buf_adj_8951[3]), .\SLO_buf[4] (SLO_buf_adj_8951[4]), 
            .\SLO_buf[5] (SLO_buf_adj_8951[5]), .\SLO_buf[6] (SLO_buf_adj_8951[6]), 
            .\SLO_buf[7] (SLO_buf_adj_8951[7]), .\SLO_buf[8] (SLO_buf_adj_8951[8]), 
            .\SLO_buf[9] (SLO_buf_adj_8951[9]), .\SLO_buf[10] (SLO_buf_adj_8951[10]), 
            .\SLO_buf[11] (SLO_buf_adj_8951[11]), .\SLO_buf[12] (SLO_buf_adj_8951[12]), 
            .\SLO_buf[13] (SLO_buf_adj_8951[13]), .\SLO_buf[14] (SLO_buf_adj_8951[14]), 
            .\SLO_buf[15] (SLO_buf_adj_8951[15]), .\SLO_buf[16] (SLO_buf_adj_8951[16]), 
            .\SLO_buf[17] (SLO_buf_adj_8951[17]), .\SLO_buf[18] (SLO_buf_adj_8951[18]), 
            .\SLO_buf[19] (SLO_buf_adj_8951[19]), .\SLO_buf[20] (SLO_buf_adj_8951[20]), 
            .\SLO_buf[21] (SLO_buf_adj_8951[21]), .\SLO_buf[22] (SLO_buf_adj_8951[22]), 
            .\SLO_buf[23] (SLO_buf_adj_8951[23]), .\SLO_buf[24] (SLO_buf_adj_8951[24]), 
            .\SLO_buf[25] (SLO_buf_adj_8951[25]), .\SLO_buf[26] (SLO_buf_adj_8951[26]), 
            .\SLO_buf[27] (SLO_buf_adj_8951[27]), .\SLO_buf[28] (SLO_buf_adj_8951[28]), 
            .\SLO_buf[29] (SLO_buf_adj_8951[29]), .\spi_data_out_r_39__N_5513[16] (spi_data_out_r_39__N_5513[16]), 
            .\spi_data_out_r_39__N_6114[1] (spi_data_out_r_39__N_6114[1]), 
            .\spi_data_out_r_39__N_5852[2] (spi_data_out_r_39__N_5852[2]), 
            .\spi_data_out_r_39__N_6114[2] (spi_data_out_r_39__N_6114[2]), 
            .\spi_data_out_r_39__N_6114[3] (spi_data_out_r_39__N_6114[3]), 
            .\spi_data_out_r_39__N_6114[4] (spi_data_out_r_39__N_6114[4]), 
            .\spi_data_out_r_39__N_6114[5] (spi_data_out_r_39__N_6114[5]), 
            .\spi_data_out_r_39__N_6114[6] (spi_data_out_r_39__N_6114[6]), 
            .\spi_data_out_r_39__N_6114[7] (spi_data_out_r_39__N_6114[7]), 
            .\spi_data_out_r_39__N_6114[8] (spi_data_out_r_39__N_6114[8]), 
            .\spi_data_out_r_39__N_6114[9] (spi_data_out_r_39__N_6114[9]), 
            .\spi_data_out_r_39__N_6114[10] (spi_data_out_r_39__N_6114[10]), 
            .\spi_data_out_r_39__N_6114[11] (spi_data_out_r_39__N_6114[11]), 
            .\spi_data_out_r_39__N_6114[12] (spi_data_out_r_39__N_6114[12]), 
            .\spi_data_out_r_39__N_6114[13] (spi_data_out_r_39__N_6114[13]), 
            .\spi_data_out_r_39__N_6114[14] (spi_data_out_r_39__N_6114[14]), 
            .\spi_data_out_r_39__N_6114[15] (spi_data_out_r_39__N_6114[15]), 
            .n29076(n29076), .\spi_data_out_r_39__N_6114[32] (spi_data_out_r_39__N_6114[32]), 
            .\spi_data_out_r_39__N_6114[33] (spi_data_out_r_39__N_6114[33]), 
            .\spi_data_out_r_39__N_6114[34] (spi_data_out_r_39__N_6114[34]), 
            .\spi_data_out_r_39__N_6114[35] (spi_data_out_r_39__N_6114[35]), 
            .\spi_data_out_r_39__N_4496[16] (spi_data_out_r_39__N_4496[16]), 
            .\spi_data_out_r_39__N_2338[2] (spi_data_out_r_39__N_2338[2]), 
            .n8(n8), .\spi_data_out_r_39__N_2998[2] (spi_data_out_r_39__N_2998[2]), 
            .clear_intrpt_adj_172(clear_intrpt_adj_7962), .n15(n15), .\spi_data_out_r_39__N_2714[2] (spi_data_out_r_39__N_2714[2]), 
            .clear_intrpt_adj_173(clear_intrpt_adj_7958), .n11(n11), .\spi_data_out_r_39__N_4835[2] (spi_data_out_r_39__N_4835[2]), 
            .n19(n19), .\spi_data_out_r_39__N_3818[16] (spi_data_out_r_39__N_3818[16]), 
            .\spi_data_out_r_39__N_4157[0] (spi_data_out_r_39__N_4157[0]), 
            .n17(n17), .\spi_data_out_r_39__N_1168[0] (spi_data_out_r_39__N_1168[0]), 
            .n3(n3_adj_8181), .\spi_data_out_r_39__N_5174[0] (spi_data_out_r_39__N_5174[0]), 
            .n20(n20), .\spi_data_out_r_39__N_2998[0] (spi_data_out_r_39__N_2998[0]), 
            .n15_adj_174(n15_adj_8184), .\spi_data_out_r_39__N_934[0] (spi_data_out_r_39__N_934[0]), 
            .n2(n2_adj_8180), .\spi_data_out_r_39__N_5513[0] (spi_data_out_r_39__N_5513[0]), 
            .n21(n21), .\spi_data_out_r_39__N_1402[0] (spi_data_out_r_39__N_1402[0]), 
            .n4_adj_175(n4_adj_8182), .\spi_data_out_r_39__N_2714[0] (spi_data_out_r_39__N_2714[0]), 
            .n11_adj_176(n11_adj_8183), .\spi_data_out_r[1] (spi_data_out_r[1]), 
            .\spi_data_out_r_39__N_2643[1] (spi_data_out_r_39__N_2643[1]), 
            .\spi_data_out_r_39__N_2856[1] (spi_data_out_r_39__N_2856[1]), 
            .clear_intrpt_adj_177(clear_intrpt_adj_7956), .\spi_data_out_r_39__N_934[1] (spi_data_out_r_39__N_934[1]), 
            .\spi_data_out_r_39__N_4157[1] (spi_data_out_r_39__N_4157[1]), 
            .\spi_data_out_r_39__N_1168[1] (spi_data_out_r_39__N_1168[1]), 
            .\spi_data_out_r_39__N_2927[1] (spi_data_out_r_39__N_2927[1]), 
            .\spi_data_out_r_39__N_2785[1] (spi_data_out_r_39__N_2785[1]), 
            .clear_intrpt_adj_178(clear_intrpt_adj_7961), .clear_intrpt_adj_179(clear_intrpt_adj_7959), 
            .\spi_data_out_r_39__N_1402[1] (spi_data_out_r_39__N_1402[1]), 
            .\spi_data_out_r_39__N_5174[1] (spi_data_out_r_39__N_5174[1]), 
            .\spi_data_out_r_39__N_3818[1] (spi_data_out_r_39__N_3818[1]), 
            .\spi_data_out_r_39__N_2338[1] (spi_data_out_r_39__N_2338[1]), 
            .\spi_data_out_r_39__N_4496[21] (spi_data_out_r_39__N_4496[21]), 
            .\spi_data_out_r_39__N_4496[1] (spi_data_out_r_39__N_4496[1]), 
            .\spi_data_out_r_39__N_1870[1] (spi_data_out_r_39__N_1870[1]), 
            .\spi_data_out_r_39__N_2998[1] (spi_data_out_r_39__N_2998[1]), 
            .\spi_data_out_r_39__N_2104[1] (spi_data_out_r_39__N_2104[1]), 
            .\spi_data_out_r_39__N_2572[1] (spi_data_out_r_39__N_2572[1]), 
            .clear_intrpt_adj_180(clear_intrpt), .\spi_data_out_r_39__N_4835[1] (spi_data_out_r_39__N_4835[1]), 
            .\spi_data_out_r_39__N_5513[1] (spi_data_out_r_39__N_5513[1]), 
            .\spi_data_out_r_39__N_1636[1] (spi_data_out_r_39__N_1636[1]), 
            .\spi_data_out_r_39__N_2714[1] (spi_data_out_r_39__N_2714[1]), 
            .\spi_data_out_r[3] (spi_data_out_r[3]), .\spi_data_out_r_39__N_1168[3] (spi_data_out_r_39__N_1168[3]), 
            .\spi_data_out_r_39__N_4835[3] (spi_data_out_r_39__N_4835[3]), 
            .\spi_data_out_r_39__N_5513[3] (spi_data_out_r_39__N_5513[3]), 
            .\spi_data_out_r_39__N_4496[3] (spi_data_out_r_39__N_4496[3]), 
            .\spi_data_out_r_39__N_3818[3] (spi_data_out_r_39__N_3818[3]), 
            .\spi_data_out_r_39__N_2104[3] (spi_data_out_r_39__N_2104[3]), 
            .\spi_data_out_r_39__N_1870[3] (spi_data_out_r_39__N_1870[3]), 
            .\spi_data_out_r_39__N_1402[3] (spi_data_out_r_39__N_1402[3]), 
            .\spi_data_out_r_39__N_2338[3] (spi_data_out_r_39__N_2338[3]), 
            .\spi_data_out_r_39__N_5174[3] (spi_data_out_r_39__N_5174[3]), 
            .\spi_data_out_r_39__N_1636[3] (spi_data_out_r_39__N_1636[3]), 
            .\spi_data_out_r_39__N_934[3] (spi_data_out_r_39__N_934[3]), .\spi_data_out_r_39__N_4157[3] (spi_data_out_r_39__N_4157[3]), 
            .\spi_data_out_r[4] (spi_data_out_r[4]), .\spi_data_out_r_39__N_1168[4] (spi_data_out_r_39__N_1168[4]), 
            .\spi_data_out_r_39__N_4835[4] (spi_data_out_r_39__N_4835[4]), 
            .\spi_data_out_r_39__N_5513[4] (spi_data_out_r_39__N_5513[4]), 
            .\spi_data_out_r_39__N_4496[4] (spi_data_out_r_39__N_4496[4]), 
            .\spi_data_out_r_39__N_2104[16] (spi_data_out_r_39__N_2104[16]), 
            .\spi_data_out_r_39__N_1870[16] (spi_data_out_r_39__N_1870[16]), 
            .\spi_data_out_r_39__N_3818[4] (spi_data_out_r_39__N_3818[4]), 
            .\spi_data_out_r_39__N_2104[4] (spi_data_out_r_39__N_2104[4]), 
            .\spi_data_out_r_39__N_1870[4] (spi_data_out_r_39__N_1870[4]), 
            .\spi_data_out_r_39__N_1402[16] (spi_data_out_r_39__N_1402[16]), 
            .\spi_data_out_r_39__N_1402[4] (spi_data_out_r_39__N_1402[4]), 
            .\spi_data_out_r_39__N_2338[4] (spi_data_out_r_39__N_2338[4]), 
            .\spi_data_out_r_39__N_5174[4] (spi_data_out_r_39__N_5174[4]), 
            .\spi_data_out_r_39__N_1636[4] (spi_data_out_r_39__N_1636[4]), 
            .\spi_data_out_r_39__N_934[4] (spi_data_out_r_39__N_934[4]), .\spi_data_out_r_39__N_4157[4] (spi_data_out_r_39__N_4157[4]), 
            .\spi_data_out_r[5] (spi_data_out_r[5]), .\spi_data_out_r_39__N_1168[5] (spi_data_out_r_39__N_1168[5]), 
            .\spi_data_out_r_39__N_4835[5] (spi_data_out_r_39__N_4835[5]), 
            .\spi_data_out_r_39__N_5513[5] (spi_data_out_r_39__N_5513[5]), 
            .\spi_data_out_r_39__N_4496[5] (spi_data_out_r_39__N_4496[5]), 
            .\spi_data_out_r_39__N_3818[5] (spi_data_out_r_39__N_3818[5]), 
            .\spi_data_out_r_39__N_2104[5] (spi_data_out_r_39__N_2104[5]), 
            .\spi_data_out_r_39__N_1870[5] (spi_data_out_r_39__N_1870[5]), 
            .\spi_data_out_r_39__N_1402[5] (spi_data_out_r_39__N_1402[5]), 
            .\spi_data_out_r_39__N_2338[5] (spi_data_out_r_39__N_2338[5]), 
            .\spi_data_out_r_39__N_5174[5] (spi_data_out_r_39__N_5174[5]), 
            .\spi_data_out_r_39__N_1636[5] (spi_data_out_r_39__N_1636[5]), 
            .\spi_data_out_r_39__N_934[5] (spi_data_out_r_39__N_934[5]), .\spi_data_out_r_39__N_4157[5] (spi_data_out_r_39__N_4157[5]), 
            .\spi_data_out_r[6] (spi_data_out_r[6]), .\spi_data_out_r_39__N_1168[6] (spi_data_out_r_39__N_1168[6]), 
            .\spi_data_out_r_39__N_4835[6] (spi_data_out_r_39__N_4835[6]), 
            .\spi_data_out_r_39__N_5513[6] (spi_data_out_r_39__N_5513[6]), 
            .\spi_data_out_r_39__N_4496[6] (spi_data_out_r_39__N_4496[6]), 
            .\spi_data_out_r_39__N_3818[6] (spi_data_out_r_39__N_3818[6]), 
            .\spi_data_out_r_39__N_2104[6] (spi_data_out_r_39__N_2104[6]), 
            .\spi_data_out_r_39__N_1870[6] (spi_data_out_r_39__N_1870[6]), 
            .\spi_data_out_r_39__N_1402[6] (spi_data_out_r_39__N_1402[6]), 
            .\spi_data_out_r_39__N_2338[6] (spi_data_out_r_39__N_2338[6]), 
            .\spi_data_out_r_39__N_5174[6] (spi_data_out_r_39__N_5174[6]), 
            .\spi_data_out_r_39__N_1636[6] (spi_data_out_r_39__N_1636[6]), 
            .\spi_data_out_r_39__N_934[6] (spi_data_out_r_39__N_934[6]), .\spi_data_out_r_39__N_4157[6] (spi_data_out_r_39__N_4157[6]), 
            .\spi_data_out_r[7] (spi_data_out_r[7]), .\spi_data_out_r_39__N_1168[7] (spi_data_out_r_39__N_1168[7]), 
            .\spi_data_out_r_39__N_4835[7] (spi_data_out_r_39__N_4835[7]), 
            .\spi_data_out_r_39__N_5513[7] (spi_data_out_r_39__N_5513[7]), 
            .\spi_data_out_r_39__N_4496[7] (spi_data_out_r_39__N_4496[7]), 
            .\spi_data_out_r_39__N_3818[7] (spi_data_out_r_39__N_3818[7]), 
            .\spi_data_out_r_39__N_2104[7] (spi_data_out_r_39__N_2104[7]), 
            .\spi_data_out_r_39__N_1870[7] (spi_data_out_r_39__N_1870[7]), 
            .\spi_data_out_r_39__N_1402[7] (spi_data_out_r_39__N_1402[7]), 
            .\spi_data_out_r_39__N_2338[7] (spi_data_out_r_39__N_2338[7]), 
            .\spi_data_out_r_39__N_5174[7] (spi_data_out_r_39__N_5174[7]), 
            .\spi_data_out_r_39__N_1636[7] (spi_data_out_r_39__N_1636[7]), 
            .\spi_data_out_r_39__N_934[7] (spi_data_out_r_39__N_934[7]), .\spi_data_out_r_39__N_4157[7] (spi_data_out_r_39__N_4157[7]), 
            .\spi_data_out_r[8] (spi_data_out_r[8]), .\spi_data_out_r_39__N_1168[8] (spi_data_out_r_39__N_1168[8]), 
            .\spi_data_out_r_39__N_4835[8] (spi_data_out_r_39__N_4835[8]), 
            .\spi_data_out_r_39__N_5513[8] (spi_data_out_r_39__N_5513[8]), 
            .\spi_data_out_r_39__N_4496[8] (spi_data_out_r_39__N_4496[8]), 
            .\spi_data_out_r_39__N_3818[8] (spi_data_out_r_39__N_3818[8]), 
            .\spi_data_out_r_39__N_2104[8] (spi_data_out_r_39__N_2104[8]), 
            .\spi_data_out_r_39__N_1870[8] (spi_data_out_r_39__N_1870[8]), 
            .\spi_data_out_r_39__N_1402[8] (spi_data_out_r_39__N_1402[8]), 
            .\spi_data_out_r_39__N_2338[8] (spi_data_out_r_39__N_2338[8]), 
            .\spi_data_out_r_39__N_5174[8] (spi_data_out_r_39__N_5174[8]), 
            .\spi_data_out_r_39__N_1636[8] (spi_data_out_r_39__N_1636[8]), 
            .\spi_data_out_r_39__N_934[8] (spi_data_out_r_39__N_934[8]), .\spi_data_out_r_39__N_4157[8] (spi_data_out_r_39__N_4157[8]), 
            .\spi_data_out_r[9] (spi_data_out_r[9]), .\spi_data_out_r_39__N_1168[9] (spi_data_out_r_39__N_1168[9]), 
            .\spi_data_out_r_39__N_4835[9] (spi_data_out_r_39__N_4835[9]), 
            .\spi_data_out_r_39__N_5513[9] (spi_data_out_r_39__N_5513[9]), 
            .\spi_data_out_r_39__N_4496[9] (spi_data_out_r_39__N_4496[9]), 
            .\spi_data_out_r_39__N_3818[9] (spi_data_out_r_39__N_3818[9]), 
            .\spi_data_out_r_39__N_2104[9] (spi_data_out_r_39__N_2104[9]), 
            .\spi_data_out_r_39__N_1870[9] (spi_data_out_r_39__N_1870[9]), 
            .\spi_data_out_r_39__N_1402[9] (spi_data_out_r_39__N_1402[9]), 
            .\spi_data_out_r_39__N_2338[9] (spi_data_out_r_39__N_2338[9]), 
            .\spi_data_out_r_39__N_5174[9] (spi_data_out_r_39__N_5174[9]), 
            .\spi_data_out_r_39__N_1636[9] (spi_data_out_r_39__N_1636[9]), 
            .\spi_data_out_r_39__N_2338[16] (spi_data_out_r_39__N_2338[16]), 
            .\spi_data_out_r_39__N_5174[16] (spi_data_out_r_39__N_5174[16]), 
            .\spi_data_out_r_39__N_934[9] (spi_data_out_r_39__N_934[9]), .\spi_data_out_r_39__N_4157[9] (spi_data_out_r_39__N_4157[9]), 
            .\spi_data_out_r[10] (spi_data_out_r[10]), .\spi_data_out_r_39__N_1168[10] (spi_data_out_r_39__N_1168[10]), 
            .\spi_data_out_r_39__N_4835[10] (spi_data_out_r_39__N_4835[10]), 
            .\spi_data_out_r_39__N_5513[10] (spi_data_out_r_39__N_5513[10]), 
            .\spi_data_out_r_39__N_4496[10] (spi_data_out_r_39__N_4496[10]), 
            .\spi_data_out_r_39__N_3818[10] (spi_data_out_r_39__N_3818[10]), 
            .\spi_data_out_r_39__N_2104[10] (spi_data_out_r_39__N_2104[10]), 
            .\spi_data_out_r_39__N_1870[10] (spi_data_out_r_39__N_1870[10]), 
            .\spi_data_out_r_39__N_1402[10] (spi_data_out_r_39__N_1402[10]), 
            .\spi_data_out_r_39__N_2338[10] (spi_data_out_r_39__N_2338[10]), 
            .\spi_data_out_r_39__N_5174[10] (spi_data_out_r_39__N_5174[10]), 
            .\spi_data_out_r_39__N_1636[10] (spi_data_out_r_39__N_1636[10]), 
            .\spi_data_out_r_39__N_934[10] (spi_data_out_r_39__N_934[10]), 
            .\spi_data_out_r_39__N_4157[10] (spi_data_out_r_39__N_4157[10]), 
            .\spi_data_out_r[11] (spi_data_out_r[11]), .\spi_data_out_r_39__N_1168[11] (spi_data_out_r_39__N_1168[11]), 
            .\spi_data_out_r_39__N_4835[11] (spi_data_out_r_39__N_4835[11]), 
            .\spi_data_out_r_39__N_5513[11] (spi_data_out_r_39__N_5513[11]), 
            .\spi_data_out_r_39__N_4496[11] (spi_data_out_r_39__N_4496[11]), 
            .\spi_data_out_r_39__N_3818[11] (spi_data_out_r_39__N_3818[11]), 
            .\spi_data_out_r_39__N_2104[11] (spi_data_out_r_39__N_2104[11]), 
            .\spi_data_out_r_39__N_1870[11] (spi_data_out_r_39__N_1870[11]), 
            .\spi_data_out_r_39__N_1402[11] (spi_data_out_r_39__N_1402[11]), 
            .\spi_data_out_r_39__N_2338[11] (spi_data_out_r_39__N_2338[11]), 
            .\spi_data_out_r_39__N_5174[11] (spi_data_out_r_39__N_5174[11]), 
            .\spi_data_out_r_39__N_1636[11] (spi_data_out_r_39__N_1636[11]), 
            .\spi_data_out_r_39__N_934[11] (spi_data_out_r_39__N_934[11]), 
            .\spi_data_out_r_39__N_4157[11] (spi_data_out_r_39__N_4157[11]), 
            .\spi_data_out_r[12] (spi_data_out_r[12]), .\spi_data_out_r_39__N_1168[12] (spi_data_out_r_39__N_1168[12]), 
            .\spi_data_out_r_39__N_4835[12] (spi_data_out_r_39__N_4835[12]), 
            .\spi_data_out_r_39__N_5513[12] (spi_data_out_r_39__N_5513[12]), 
            .\spi_data_out_r_39__N_4496[12] (spi_data_out_r_39__N_4496[12]), 
            .\spi_data_out_r_39__N_3818[12] (spi_data_out_r_39__N_3818[12]), 
            .\spi_data_out_r_39__N_2104[12] (spi_data_out_r_39__N_2104[12]), 
            .\spi_data_out_r_39__N_1870[12] (spi_data_out_r_39__N_1870[12]), 
            .\spi_data_out_r_39__N_1402[12] (spi_data_out_r_39__N_1402[12]), 
            .\spi_data_out_r_39__N_2338[12] (spi_data_out_r_39__N_2338[12]), 
            .\spi_data_out_r_39__N_5174[12] (spi_data_out_r_39__N_5174[12]), 
            .\spi_data_out_r_39__N_1636[12] (spi_data_out_r_39__N_1636[12]), 
            .\spi_data_out_r_39__N_934[12] (spi_data_out_r_39__N_934[12]), 
            .\spi_data_out_r_39__N_4157[12] (spi_data_out_r_39__N_4157[12]), 
            .\spi_data_out_r[13] (spi_data_out_r[13]), .\spi_data_out_r_39__N_1168[13] (spi_data_out_r_39__N_1168[13]), 
            .\spi_data_out_r_39__N_4835[13] (spi_data_out_r_39__N_4835[13]), 
            .\spi_data_out_r_39__N_5513[13] (spi_data_out_r_39__N_5513[13]), 
            .\spi_data_out_r_39__N_4496[13] (spi_data_out_r_39__N_4496[13]), 
            .\spi_data_out_r_39__N_3818[13] (spi_data_out_r_39__N_3818[13]), 
            .\spi_data_out_r_39__N_2104[13] (spi_data_out_r_39__N_2104[13]), 
            .\spi_data_out_r_39__N_1870[13] (spi_data_out_r_39__N_1870[13]), 
            .\spi_data_out_r_39__N_1402[13] (spi_data_out_r_39__N_1402[13]), 
            .\spi_data_out_r_39__N_2338[13] (spi_data_out_r_39__N_2338[13]), 
            .\spi_data_out_r_39__N_5174[13] (spi_data_out_r_39__N_5174[13]), 
            .\spi_data_out_r_39__N_1636[13] (spi_data_out_r_39__N_1636[13]), 
            .\spi_data_out_r_39__N_934[13] (spi_data_out_r_39__N_934[13]), 
            .\spi_data_out_r_39__N_4157[13] (spi_data_out_r_39__N_4157[13]), 
            .\spi_data_out_r[14] (spi_data_out_r[14]), .\spi_data_out_r_39__N_1168[14] (spi_data_out_r_39__N_1168[14]), 
            .\spi_data_out_r_39__N_4835[14] (spi_data_out_r_39__N_4835[14]), 
            .\spi_data_out_r_39__N_5513[14] (spi_data_out_r_39__N_5513[14]), 
            .\spi_data_out_r_39__N_4496[14] (spi_data_out_r_39__N_4496[14]), 
            .\spi_data_out_r_39__N_3818[14] (spi_data_out_r_39__N_3818[14]), 
            .\spi_data_out_r_39__N_2104[14] (spi_data_out_r_39__N_2104[14]), 
            .\spi_data_out_r_39__N_1870[14] (spi_data_out_r_39__N_1870[14]), 
            .\spi_data_out_r_39__N_1402[14] (spi_data_out_r_39__N_1402[14]), 
            .\spi_data_out_r_39__N_2338[14] (spi_data_out_r_39__N_2338[14]), 
            .\spi_data_out_r_39__N_5174[14] (spi_data_out_r_39__N_5174[14]), 
            .\spi_data_out_r_39__N_1636[14] (spi_data_out_r_39__N_1636[14]), 
            .\spi_data_out_r_39__N_934[14] (spi_data_out_r_39__N_934[14]), 
            .\spi_data_out_r_39__N_4157[14] (spi_data_out_r_39__N_4157[14]), 
            .\spi_data_out_r[15] (spi_data_out_r[15]), .\spi_data_out_r_39__N_1168[15] (spi_data_out_r_39__N_1168[15]), 
            .\spi_data_out_r_39__N_4835[15] (spi_data_out_r_39__N_4835[15]), 
            .\spi_data_out_r_39__N_1636[16] (spi_data_out_r_39__N_1636[16]), 
            .\spi_data_out_r_39__N_5513[15] (spi_data_out_r_39__N_5513[15]), 
            .\spi_data_out_r_39__N_4496[15] (spi_data_out_r_39__N_4496[15]), 
            .\spi_data_out_r_39__N_3818[15] (spi_data_out_r_39__N_3818[15]), 
            .\spi_data_out_r_39__N_2104[15] (spi_data_out_r_39__N_2104[15]), 
            .\spi_data_out_r_39__N_1870[15] (spi_data_out_r_39__N_1870[15]), 
            .\spi_data_out_r_39__N_1402[15] (spi_data_out_r_39__N_1402[15]), 
            .\spi_data_out_r_39__N_2338[15] (spi_data_out_r_39__N_2338[15]), 
            .\spi_data_out_r_39__N_5174[15] (spi_data_out_r_39__N_5174[15]), 
            .\spi_data_out_r_39__N_934[16] (spi_data_out_r_39__N_934[16]), 
            .\spi_data_out_r_39__N_4157[16] (spi_data_out_r_39__N_4157[16]), 
            .\spi_data_out_r[17] (spi_data_out_r[17]), .\spi_data_out_r_39__N_1168[17] (spi_data_out_r_39__N_1168[17]), 
            .\spi_data_out_r_39__N_4835[17] (spi_data_out_r_39__N_4835[17]), 
            .\spi_data_out_r_39__N_5513[17] (spi_data_out_r_39__N_5513[17]), 
            .\spi_data_out_r_39__N_4496[17] (spi_data_out_r_39__N_4496[17]), 
            .\spi_data_out_r_39__N_3818[17] (spi_data_out_r_39__N_3818[17]), 
            .\spi_data_out_r_39__N_2104[17] (spi_data_out_r_39__N_2104[17]), 
            .\spi_data_out_r_39__N_1870[17] (spi_data_out_r_39__N_1870[17]), 
            .\spi_data_out_r_39__N_1402[17] (spi_data_out_r_39__N_1402[17]), 
            .\spi_data_out_r_39__N_2338[17] (spi_data_out_r_39__N_2338[17]), 
            .\spi_data_out_r_39__N_5174[17] (spi_data_out_r_39__N_5174[17]), 
            .\spi_data_out_r_39__N_1636[17] (spi_data_out_r_39__N_1636[17]), 
            .\spi_data_out_r_39__N_934[17] (spi_data_out_r_39__N_934[17]), 
            .\spi_data_out_r_39__N_4157[17] (spi_data_out_r_39__N_4157[17]), 
            .\spi_data_out_r[18] (spi_data_out_r[18]), .\spi_data_out_r_39__N_1168[18] (spi_data_out_r_39__N_1168[18]), 
            .\spi_data_out_r_39__N_4835[18] (spi_data_out_r_39__N_4835[18]), 
            .\spi_data_out_r_39__N_5513[18] (spi_data_out_r_39__N_5513[18]), 
            .\spi_data_out_r_39__N_4496[18] (spi_data_out_r_39__N_4496[18]), 
            .\spi_data_out_r_39__N_3818[18] (spi_data_out_r_39__N_3818[18]), 
            .\spi_data_out_r_39__N_2104[18] (spi_data_out_r_39__N_2104[18]), 
            .\spi_data_out_r_39__N_1870[18] (spi_data_out_r_39__N_1870[18]), 
            .\spi_data_out_r_39__N_1402[18] (spi_data_out_r_39__N_1402[18]), 
            .\spi_data_out_r_39__N_2338[18] (spi_data_out_r_39__N_2338[18]), 
            .\spi_data_out_r_39__N_5174[18] (spi_data_out_r_39__N_5174[18]), 
            .\spi_data_out_r_39__N_1636[18] (spi_data_out_r_39__N_1636[18]), 
            .\spi_data_out_r_39__N_934[18] (spi_data_out_r_39__N_934[18]), 
            .\spi_data_out_r_39__N_4157[18] (spi_data_out_r_39__N_4157[18]), 
            .\spi_data_out_r[19] (spi_data_out_r[19]), .\spi_data_out_r_39__N_1168[19] (spi_data_out_r_39__N_1168[19]), 
            .\spi_data_out_r_39__N_4835[19] (spi_data_out_r_39__N_4835[19]), 
            .\spi_data_out_r_39__N_5513[19] (spi_data_out_r_39__N_5513[19]), 
            .\spi_data_out_r_39__N_4496[19] (spi_data_out_r_39__N_4496[19]), 
            .\spi_data_out_r_39__N_3818[19] (spi_data_out_r_39__N_3818[19]), 
            .\spi_data_out_r_39__N_2104[19] (spi_data_out_r_39__N_2104[19]), 
            .\spi_data_out_r_39__N_1870[19] (spi_data_out_r_39__N_1870[19]), 
            .\spi_data_out_r_39__N_1402[19] (spi_data_out_r_39__N_1402[19]), 
            .\spi_data_out_r_39__N_2338[19] (spi_data_out_r_39__N_2338[19]), 
            .\spi_data_out_r_39__N_5174[19] (spi_data_out_r_39__N_5174[19]), 
            .\spi_data_out_r_39__N_1636[19] (spi_data_out_r_39__N_1636[19]), 
            .\spi_data_out_r_39__N_934[19] (spi_data_out_r_39__N_934[19]), 
            .\spi_data_out_r_39__N_4157[19] (spi_data_out_r_39__N_4157[19]), 
            .\spi_data_out_r[20] (spi_data_out_r[20]), .\spi_data_out_r_39__N_1168[20] (spi_data_out_r_39__N_1168[20]), 
            .reset_r(reset_r_adj_8089), .clk_enable_521(clk_enable_521), 
            .n29083(n29083), .\spi_data_out_r_39__N_4835[20] (spi_data_out_r_39__N_4835[20]), 
            .\spi_data_out_r_39__N_5513[20] (spi_data_out_r_39__N_5513[20]), 
            .\spi_data_out_r_39__N_4496[20] (spi_data_out_r_39__N_4496[20]), 
            .\spi_data_out_r_39__N_3818[20] (spi_data_out_r_39__N_3818[20]), 
            .\spi_data_out_r_39__N_2104[20] (spi_data_out_r_39__N_2104[20]), 
            .\spi_data_out_r_39__N_1870[20] (spi_data_out_r_39__N_1870[20]), 
            .\spi_data_out_r_39__N_1402[20] (spi_data_out_r_39__N_1402[20]), 
            .\spi_data_out_r_39__N_2338[20] (spi_data_out_r_39__N_2338[20]), 
            .\spi_data_out_r_39__N_5174[20] (spi_data_out_r_39__N_5174[20]), 
            .\spi_data_out_r_39__N_1636[20] (spi_data_out_r_39__N_1636[20]), 
            .\spi_data_out_r_39__N_934[20] (spi_data_out_r_39__N_934[20]), 
            .\spi_data_out_r_39__N_4157[20] (spi_data_out_r_39__N_4157[20]), 
            .\spi_data_out_r[21] (spi_data_out_r[21]), .\spi_data_out_r_39__N_1168[21] (spi_data_out_r_39__N_1168[21]), 
            .\spi_data_out_r_39__N_3818[21] (spi_data_out_r_39__N_3818[21]), 
            .\spi_data_out_r_39__N_2104[21] (spi_data_out_r_39__N_2104[21]), 
            .\spi_data_out_r_39__N_1870[21] (spi_data_out_r_39__N_1870[21]), 
            .\spi_data_out_r_39__N_1402[21] (spi_data_out_r_39__N_1402[21]), 
            .\spi_data_out_r_39__N_2338[21] (spi_data_out_r_39__N_2338[21]), 
            .\spi_data_out_r_39__N_5174[21] (spi_data_out_r_39__N_5174[21])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(364[3] 407[2])
    spi_slave_top spi_slave_top_inst (.spi_addr_r({Open_0, Open_1, Open_2, 
            Open_3, Open_4, Open_5, Open_6, spi_addr_r[0]}), .clk(clk), 
            .n29247(n29247), .spi_addr({Open_7, Open_8, Open_9, Open_10, 
            Open_11, Open_12, Open_13, spi_addr[0]}), .n29239(n29239), 
            .\spi_addr_r[3] (spi_addr_r[3]), .\spi_addr[3] (spi_addr[3]), 
            .\spi_addr_r[2] (spi_addr_r[2]), .\spi_addr[2] (spi_addr[2]), 
            .\spi_addr_r[1] (spi_addr_r[1]), .\spi_addr[1] (spi_addr[1]), 
            .spi_cmd_r({Open_14, Open_15, Open_16, Open_17, Open_18, 
            Open_19, Open_20, Open_21, Open_22, Open_23, Open_24, 
            Open_25, spi_cmd_r[3:0]}), .\spi_data_r[0] (spi_data_r[0]), 
            .clk_enable_524(clk_enable_524), .n27(n27), .n29182(n29182), 
            .n13074(n13074), .n29077(n29077), .n29761(n29761), .n27256(n27256), 
            .n29174(n29174), .n29211(n29211), .spi_addr_valid(spi_addr_valid), 
            .spi_cmd_valid(spi_cmd_valid), .resetn_c(resetn_c), .spi_scsn_c(spi_scsn_c), 
            .spi_sdo_valid_N_296(spi_sdo_valid_N_296), .n29162(n29162), 
            .n29161(n29161), .n29144(n29144), .n29122(n29122), .n29251(n29251), 
            .n29254(n29254), .n27283(n27283), .n29216(n29216), .n27058(n27058), 
            .n29169(n29169), .n6(n6), .n13265(n13265), .n29214(n29214), 
            .n29127(n29127), .n29118(n29118), .n29130(n29130), .\spi_data_r[31] (spi_data_r[31]), 
            .\spi_data_r[30] (spi_data_r[30]), .\spi_data_r[29] (spi_data_r[29]), 
            .\spi_data_r[28] (spi_data_r[28]), .\spi_data_r[27] (spi_data_r[27]), 
            .\spi_data_r[26] (spi_data_r[26]), .\spi_data_r[25] (spi_data_r[25]), 
            .\spi_data_r[24] (spi_data_r[24]), .\spi_data_r[23] (spi_data_r[23]), 
            .\spi_data_r[22] (spi_data_r[22]), .\spi_data_r[21] (spi_data_r[21]), 
            .\spi_data_r[20] (spi_data_r[20]), .\spi_data_r[19] (spi_data_r[19]), 
            .\spi_data_r[18] (spi_data_r[18]), .\spi_data_r[17] (spi_data_r[17]), 
            .\spi_data_r[16] (spi_data_r[16]), .\spi_data_r[15] (spi_data_r[15]), 
            .\spi_data_r[14] (spi_data_r[14]), .\spi_data_r[13] (spi_data_r[13]), 
            .\spi_data_r[12] (spi_data_r[12]), .\spi_data_r[11] (spi_data_r[11]), 
            .\spi_data_r[10] (spi_data_r[10]), .\spi_data_r[9] (spi_data_r[9]), 
            .\spi_data_r[8] (spi_data_r[8]), .\spi_data_r[7] (spi_data_r[7]), 
            .\spi_data_r[6] (spi_data_r[6]), .\spi_data_r[5] (spi_data_r[5]), 
            .\spi_data_r[4] (spi_data_r[4]), .\spi_data_r[3] (spi_data_r[3]), 
            .\spi_data_r[2] (spi_data_r[2]), .\spi_data_r[1] (spi_data_r[1]), 
            .n27338(n27338), .n29311(n29311), .n27259(n27259), .n29287(n29287), 
            .n29255(n29255), .reset_r_N_4813(reset_r_N_4813), .clk_enable_190(clk_enable_190), 
            .n65(n65_adj_8152), .n29070(n29070), .spi_sdo_valid_N_297(spi_sdo_valid_N_297), 
            .\spi_data_out_r_39__N_2643[2] (spi_data_out_r_39__N_2643[2]), 
            .n13(n13), .clear_intrpt(clear_intrpt_adj_7956), .n4(n4), 
            .\spi_data_out_r_39__N_934[2] (spi_data_out_r_39__N_934[2]), .n19(n19), 
            .spi_data_out_r_39__N_974(spi_data_out_r_39__N_974), .spi_data_valid_r(spi_data_valid_r), 
            .spi_data_valid(spi_data_valid), .spi_cmd({Open_26, Open_27, 
            Open_28, Open_29, Open_30, Open_31, Open_32, Open_33, 
            Open_34, Open_35, Open_36, Open_37, Open_38, spi_cmd[2:1], 
            Open_39}), .\spi_data_out_r_39__N_4157[2] (spi_data_out_r_39__N_4157[2]), 
            .\spi_data_out_r_39__N_1168[2] (spi_data_out_r_39__N_1168[2]), 
            .spi_data_out_r_39__N_4197(spi_data_out_r_39__N_4197), .spi_data_out_r_39__N_1208(spi_data_out_r_39__N_1208), 
            .\spi_data_out_r_39__N_2927[2] (spi_data_out_r_39__N_2927[2]), 
            .\spi_data_out_r_39__N_2785[2] (spi_data_out_r_39__N_2785[2]), 
            .clear_intrpt_adj_151(clear_intrpt_adj_7961), .clear_intrpt_adj_152(clear_intrpt_adj_7959), 
            .n8(n8), .n15(n15), .\spi_cmd[4] (spi_cmd[4]), .\spi_cmd_r[6] (spi_cmd_r[6]), 
            .\spi_cmd_r[7] (spi_cmd_r[7]), .\spi_cmd_r[8] (spi_cmd_r[8]), 
            .\spi_cmd_r[9] (spi_cmd_r[9]), .\spi_cmd_r[10] (spi_cmd_r[10]), 
            .\spi_cmd_r[11] (spi_cmd_r[11]), .\spi_cmd_r[12] (spi_cmd_r[12]), 
            .\spi_cmd_r[13] (spi_cmd_r[13]), .\spi_cmd_r[14] (spi_cmd_r[14]), 
            .\spi_cmd_r[15] (spi_cmd_r[15]), .\spi_cmd[15] (spi_cmd[15]), 
            .\spi_data_out_r[1] (spi_data_out_r[1]), .\spi_data_out_r[3] (spi_data_out_r[3]), 
            .\spi_data_out_r[4] (spi_data_out_r[4]), .\spi_data_out_r[5] (spi_data_out_r[5]), 
            .\spi_data_out_r[6] (spi_data_out_r[6]), .\spi_data_out_r[7] (spi_data_out_r[7]), 
            .\spi_data_out_r[8] (spi_data_out_r[8]), .\spi_data_out_r[9] (spi_data_out_r[9]), 
            .\spi_data_out_r[10] (spi_data_out_r[10]), .\spi_data_out_r[11] (spi_data_out_r[11]), 
            .\spi_data_out_r[12] (spi_data_out_r[12]), .\spi_data_out_r[13] (spi_data_out_r[13]), 
            .\spi_data_out_r[14] (spi_data_out_r[14]), .\spi_data_out_r[15] (spi_data_out_r[15]), 
            .\spi_data_out_r[16] (spi_data_out_r[16]), .\spi_data_out_r[17] (spi_data_out_r[17]), 
            .\spi_data_out_r[18] (spi_data_out_r[18]), .\spi_data_out_r[19] (spi_data_out_r[19]), 
            .\spi_data_out_r[20] (spi_data_out_r[20]), .\spi_data_out_r[21] (spi_data_out_r[21]), 
            .\spi_data_out_r[22] (spi_data_out_r[22]), .\spi_data_out_r[23] (spi_data_out_r[23]), 
            .\spi_data_out_r[24] (spi_data_out_r[24]), .\spi_data_out_r[25] (spi_data_out_r[25]), 
            .\spi_data_out_r[26] (spi_data_out_r[26]), .\spi_data_out_r[27] (spi_data_out_r[27]), 
            .\spi_data_out_r[28] (spi_data_out_r[28]), .\spi_data_out_r[29] (spi_data_out_r[29]), 
            .\spi_data_out_r[30] (spi_data_out_r[30]), .\spi_data_out_r[31] (spi_data_out_r[31]), 
            .\spi_data_out_r[32] (spi_data_out_r[32]), .\spi_data_out_r[33] (spi_data_out_r[33]), 
            .\spi_data_out_r[34] (spi_data_out_r[34]), .\spi_data_out_r[35] (spi_data_out_r[35]), 
            .\spi_data_out_r[36] (spi_data_out_r[36]), .\spi_data_out_r[37] (spi_data_out_r[37]), 
            .\spi_data_out_r[38] (spi_data_out_r[38]), .\spi_data_out_r[39] (spi_data_out_r[39]), 
            .\spi_data_out_r_39__N_5174[2] (spi_data_out_r_39__N_5174[2]), 
            .\spi_data_out_r_39__N_3818[2] (spi_data_out_r_39__N_3818[2]), 
            .spi_data_out_r_39__N_5214(spi_data_out_r_39__N_5214), .spi_data_out_r_39__N_3858(spi_data_out_r_39__N_3858), 
            .\spi_data_out_r_39__N_5852[2] (spi_data_out_r_39__N_5852[2]), 
            .n11(n11), .spi_data_out_r_39__N_5892(spi_data_out_r_39__N_5892), 
            .\spi_data_out_r_39__N_4496[2] (spi_data_out_r_39__N_4496[2]), 
            .\spi_data_out_r_39__N_1870[2] (spi_data_out_r_39__N_1870[2]), 
            .spi_data_out_r_39__N_4536(spi_data_out_r_39__N_4536), .spi_data_out_r_39__N_1910(spi_data_out_r_39__N_1910), 
            .\spi_data_out_r_39__N_5513[2] (spi_data_out_r_39__N_5513[2]), 
            .\spi_data_out_r_39__N_1636[2] (spi_data_out_r_39__N_1636[2]), 
            .spi_data_out_r_39__N_5553(spi_data_out_r_39__N_5553), .spi_data_out_r_39__N_1676(spi_data_out_r_39__N_1676), 
            .\spi_data_out_r_39__N_2104[2] (spi_data_out_r_39__N_2104[2]), 
            .\spi_data_out_r_39__N_2572[2] (spi_data_out_r_39__N_2572[2]), 
            .spi_data_out_r_39__N_2144(spi_data_out_r_39__N_2144), .clear_intrpt_adj_153(clear_intrpt), 
            .n29075(n29075), .n29078(n29078), .n29079(n29079), .n29080(n29080), 
            .n27286(n27286), .n65_adj_154(n65), .n29092(n29092), .\spi_data_out_r_39__N_2927[0] (spi_data_out_r_39__N_2927[0]), 
            .n17(n17), .n3(n3_adj_8181), .n20(n20), .\spi_data_out_r_39__N_3818[0] (spi_data_out_r_39__N_3818[0]), 
            .n4_adj_155(n4_adj_8182), .\spi_data_out_r_39__N_1870[0] (spi_data_out_r_39__N_1870[0]), 
            .\spi_data_out_r_39__N_2785[0] (spi_data_out_r_39__N_2785[0]), 
            .n15_adj_156(n15_adj_8184), .n2(n2_adj_8180), .\spi_data_out_r_39__N_4496[0] (spi_data_out_r_39__N_4496[0]), 
            .n11_adj_157(n11_adj_8183), .\spi_data_out_r_39__N_4835[0] (spi_data_out_r_39__N_4835[0]), 
            .n21(n21), .spi_data_out_r_39__N_4875(spi_data_out_r_39__N_4875), 
            .\spi_data_out_r_39__N_770[0] (spi_data_out_r_39__N_770[0]), .\spi_data_out_r_39__N_5852[0] (spi_data_out_r_39__N_5852[0]), 
            .spi_data_out_r_39__N_810(spi_data_out_r_39__N_810), .\spi_data_out_r_39__N_2338[0] (spi_data_out_r_39__N_2338[0]), 
            .\spi_data_out_r_39__N_2572[0] (spi_data_out_r_39__N_2572[0]), 
            .spi_data_out_r_39__N_2378(spi_data_out_r_39__N_2378), .\spi_data_out_r_39__N_2104[0] (spi_data_out_r_39__N_2104[0]), 
            .\spi_data_out_r_39__N_2856[0] (spi_data_out_r_39__N_2856[0]), 
            .clear_intrpt_adj_158(clear_intrpt_adj_7960), .\spi_data_out_r_39__N_1636[0] (spi_data_out_r_39__N_1636[0]), 
            .\spi_data_out_r_39__N_2643[0] (spi_data_out_r_39__N_2643[0]), 
            .n29089(n29089), .clk_enable_206(clk_enable_206), .n29096(n29096), 
            .n29213(n29213), .n29097(n29097), .n29106(n29106), .n29123(n29123), 
            .n29762(n29762), .n29757(n29757), .GND_net(GND_net), .spi_mosi_oe(spi_mosi_oe), 
            .spi_mosi_o(spi_mosi_o), .spi_miso_oe(spi_miso_oe), .spi_miso_o(spi_miso_o), 
            .spi_clk_oe(spi_clk_oe), .spi_clk_o(spi_clk_o), .spi_mosi_i(spi_mosi_i), 
            .spi_miso_i(spi_miso_i), .spi_clk_i(spi_clk_i), .VCC_net(VCC_net), 
            .mem_rdata_update_N_729(mem_rdata_update_N_729), .quad_set_complete(quad_set_complete_adj_7757), 
            .clk_enable_518(clk_enable_518), .n27225(n27225), .clk_enable_398(clk_enable_398), 
            .n29102(n29102), .clk_enable_188(clk_enable_188), .clk_enable_303(clk_enable_303), 
            .n32(n32), .\quad_homing[1] (quad_homing_adj_8461[1]), .n27657(n27657), 
            .n24(n24), .clk_enable_179(clk_enable_179), .clk_enable_182(clk_enable_182), 
            .intrpt_out_N_2848(intrpt_out_N_2848), .n29100(n29100), .clk_enable_185(clk_enable_185), 
            .n29134(n29134), .clk_enable_509(clk_enable_509), .EM_STOP(EM_STOP), 
            .clk_enable_306(clk_enable_306), .n29101(n29101), .clk_enable_186(clk_enable_186), 
            .quad_set_complete_adj_159(quad_set_complete_adj_7689), .n29120(n29120), 
            .clk_enable_505(clk_enable_505), .clk_enable_76(clk_enable_76), 
            .n29104(n29104), .clk_enable_436(clk_enable_436), .n19233(n19233), 
            .clk_enable_184(clk_enable_184), .clk_enable_204(clk_enable_204), 
            .intrpt_out_N_2635(intrpt_out_N_2635), .n29288(n29288), .clk_enable_183(clk_enable_183), 
            .clk_enable_271(clk_enable_271), .n29083(n29083), .clk_enable_521(clk_enable_521), 
            .quad_set_valid(quad_set_valid_adj_7824), .n66(n66), .n21446(n21446), 
            .clk_1MHz_enable_171(clk_1MHz_enable_171), .n29124(n29124), 
            .clk_enable_197(clk_enable_197), .n26948(n26948), .n13_adj_160(n13_adj_7890), 
            .n12714(n12714), .n27301(n27301), .clk_enable_193(clk_enable_193), 
            .clk_enable_200(clk_enable_200), .n29307(n29307), .clk_enable_499(clk_enable_499), 
            .n27240(n27240), .clk_enable_32(clk_enable_32), .quad_set_complete_adj_161(quad_set_complete_adj_7891), 
            .clk_enable_520(clk_enable_520), .n29286(n29286), .clk_enable_77(clk_enable_77), 
            .intrpt_out_N_2706(intrpt_out_N_2706), .quad_set_valid_adj_162(quad_set_valid), 
            .n79(n79), .n20819(n20819), .clk_1MHz_enable_340(clk_1MHz_enable_340), 
            .n27285(n27285), .n29110(n29110), .clk_enable_340(clk_enable_340), 
            .n31(n31), .\quad_homing[1]_adj_163 (quad_homing[1]), .n5(n5_adj_8136), 
            .n26(n26), .n27234(n27234), .clk_enable_174(clk_enable_174), 
            .clk_enable_171(clk_enable_171), .clk_enable_172(clk_enable_172), 
            .clk_enable_435(clk_enable_435), .n29082(n29082), .clk_enable_506(clk_enable_506), 
            .clk_enable_269(clk_enable_269), .clk_enable_167(clk_enable_167), 
            .clk_enable_28(clk_enable_28), .clk_enable_131(clk_enable_131), 
            .intrpt_out_N_2919(intrpt_out_N_2919), .clk_enable_194(clk_enable_194), 
            .clk_enable_177(clk_enable_177), .clk_enable_189(clk_enable_189), 
            .clk_enable_180(clk_enable_180), .clk_enable_162(clk_enable_162), 
            .clk_enable_166(clk_enable_166), .n29256(n29256), .clk_enable_175(clk_enable_175), 
            .clk_enable_176(clk_enable_176), .quad_set_complete_adj_164(quad_set_complete_adj_7619), 
            .n29105(n29105), .clk_enable_502(clk_enable_502), .clk_enable_526(clk_enable_526), 
            .clk_enable_342(clk_enable_342), .clk_enable_202(clk_enable_202), 
            .intrpt_out_N_2990(intrpt_out_N_2990), .clk_enable_201(clk_enable_201), 
            .clk_enable_467(clk_enable_467), .clk_enable_191(clk_enable_191), 
            .clk_enable_187(clk_enable_187), .clk_enable_192(clk_enable_192), 
            .quad_set_complete_adj_165(quad_set_complete_adj_7825), .clk_enable_519(clk_enable_519), 
            .clk_enable_170(clk_enable_170), .clk_enable_286(clk_enable_286), 
            .clk_enable_359(clk_enable_359), .reset_r_N_4474(reset_r_N_4474), 
            .clk_enable_307(clk_enable_307), .clear_intrpt_adj_166(clear_intrpt_adj_7962), 
            .intrpt_out_N_3061(intrpt_out_N_3061), .clk_enable_86(clk_enable_86), 
            .clk_enable_181(clk_enable_181), .clk_enable_288(clk_enable_288), 
            .clk_enable_433(clk_enable_433), .clk_enable_434(clk_enable_434), 
            .quad_set_complete_adj_167(quad_set_complete), .clk_enable_501(clk_enable_501), 
            .n29205(n29205), .clk_enable_169(clk_enable_169), .clear_intrpt_adj_168(clear_intrpt_adj_7958), 
            .intrpt_out_N_2777(intrpt_out_N_2777), .clk_enable_400(clk_enable_400), 
            .clk_enable_402(clk_enable_402), .quad_set_complete_adj_169(quad_set_complete_adj_7623), 
            .clk_enable_503(clk_enable_503), .clk_enable_30(clk_enable_30), 
            .n9633(n9633), .n27465(n27465), .n26928(n26928), .n29141(n29141), 
            .n29126(n29126), .n27618(n27618), .n29114(n29114), .clk_enable_20(clk_enable_20), 
            .\spi_cmd[0] (spi_cmd[0]), .n31_adj_170(n31_adj_8153)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(186[3] 206[2])
    \quad_decoder(DEV_ID=5)  \quad_ins_5..u_quad_decoder  (.quad_homing({quad_homing_adj_8461}), 
            .n29220(n29220), .pin_io_out_54(pin_io_out_54), .n95(n95), 
            .n66(n66), .n5647(n5647), .n24(n24), .n32(n32), .quad_count({quad_count_adj_8462}), 
            .clk_1MHz(clk_1MHz), .clk_1MHz_enable_171(clk_1MHz_enable_171), 
            .\spi_data_out_r_39__N_2104[0] (spi_data_out_r_39__N_2104[0]), 
            .clk(clk), .\spi_data_out_r_39__N_2249[0] (spi_data_out_r_39__N_2249[0]), 
            .\quad_b[5] (quad_b[5]), .quad_buffer({quad_buffer_adj_8463}), 
            .\mode[2]_derived_32 (mode_2_derived_32_adj_8049), .clk_enable_28(clk_enable_28), 
            .n29239(n29239), .\spi_data_r[1] (spi_data_r[1]), .n29762(n29762), 
            .clk_enable_131(clk_enable_131), .\spi_data_r[0] (spi_data_r[0]), 
            .\spi_data_r[31] (spi_data_r[31]), .\spi_data_r[30] (spi_data_r[30]), 
            .\spi_data_r[29] (spi_data_r[29]), .\spi_data_r[28] (spi_data_r[28]), 
            .\spi_data_r[27] (spi_data_r[27]), .\spi_data_r[26] (spi_data_r[26]), 
            .\spi_data_r[25] (spi_data_r[25]), .\spi_data_r[24] (spi_data_r[24]), 
            .\spi_data_r[23] (spi_data_r[23]), .\spi_data_r[22] (spi_data_r[22]), 
            .\spi_data_r[21] (spi_data_r[21]), .\spi_data_r[20] (spi_data_r[20]), 
            .\spi_data_r[19] (spi_data_r[19]), .\spi_data_r[18] (spi_data_r[18]), 
            .\spi_data_r[17] (spi_data_r[17]), .\spi_data_r[16] (spi_data_r[16]), 
            .\spi_data_r[15] (spi_data_r[15]), .\spi_data_r[14] (spi_data_r[14]), 
            .\spi_data_r[13] (spi_data_r[13]), .\spi_data_r[12] (spi_data_r[12]), 
            .\spi_data_r[11] (spi_data_r[11]), .\spi_data_r[10] (spi_data_r[10]), 
            .\spi_data_r[9] (spi_data_r[9]), .\spi_data_r[8] (spi_data_r[8]), 
            .\spi_data_r[7] (spi_data_r[7]), .\spi_data_r[6] (spi_data_r[6]), 
            .\spi_data_r[5] (spi_data_r[5]), .\spi_data_r[4] (spi_data_r[4]), 
            .\spi_data_r[3] (spi_data_r[3]), .\spi_data_r[2] (spi_data_r[2]), 
            .n29336(n29336), .spi_data_out_r_39__N_2144(spi_data_out_r_39__N_2144), 
            .spi_data_out_r_39__N_2332(spi_data_out_r_39__N_2332), .quad_set_complete(quad_set_complete_adj_7825), 
            .quad_set_valid(quad_set_valid_adj_7824), .\quad_a[5] (quad_a[5]), 
            .\spi_data_out_r_39__N_2104[31] (spi_data_out_r_39__N_2104[31]), 
            .\spi_data_out_r_39__N_2249[31] (spi_data_out_r_39__N_2249[31]), 
            .\spi_data_out_r_39__N_2104[30] (spi_data_out_r_39__N_2104[30]), 
            .\spi_data_out_r_39__N_2249[30] (spi_data_out_r_39__N_2249[30]), 
            .\spi_data_out_r_39__N_2104[29] (spi_data_out_r_39__N_2104[29]), 
            .\spi_data_out_r_39__N_2249[29] (spi_data_out_r_39__N_2249[29]), 
            .\spi_data_out_r_39__N_2104[28] (spi_data_out_r_39__N_2104[28]), 
            .\spi_data_out_r_39__N_2249[28] (spi_data_out_r_39__N_2249[28]), 
            .\spi_data_out_r_39__N_2104[27] (spi_data_out_r_39__N_2104[27]), 
            .\spi_data_out_r_39__N_2249[27] (spi_data_out_r_39__N_2249[27]), 
            .\spi_data_out_r_39__N_2104[26] (spi_data_out_r_39__N_2104[26]), 
            .\spi_data_out_r_39__N_2249[26] (spi_data_out_r_39__N_2249[26]), 
            .\spi_data_out_r_39__N_2104[25] (spi_data_out_r_39__N_2104[25]), 
            .\spi_data_out_r_39__N_2249[25] (spi_data_out_r_39__N_2249[25]), 
            .\spi_data_out_r_39__N_2104[24] (spi_data_out_r_39__N_2104[24]), 
            .\spi_data_out_r_39__N_2249[24] (spi_data_out_r_39__N_2249[24]), 
            .\spi_data_out_r_39__N_2104[23] (spi_data_out_r_39__N_2104[23]), 
            .\spi_data_out_r_39__N_2249[23] (spi_data_out_r_39__N_2249[23]), 
            .\spi_data_out_r_39__N_2104[22] (spi_data_out_r_39__N_2104[22]), 
            .\spi_data_out_r_39__N_2249[22] (spi_data_out_r_39__N_2249[22]), 
            .\spi_data_out_r_39__N_2104[21] (spi_data_out_r_39__N_2104[21]), 
            .\spi_data_out_r_39__N_2249[21] (spi_data_out_r_39__N_2249[21]), 
            .\spi_data_out_r_39__N_2104[20] (spi_data_out_r_39__N_2104[20]), 
            .\spi_data_out_r_39__N_2249[20] (spi_data_out_r_39__N_2249[20]), 
            .\spi_data_out_r_39__N_2104[19] (spi_data_out_r_39__N_2104[19]), 
            .\spi_data_out_r_39__N_2249[19] (spi_data_out_r_39__N_2249[19]), 
            .\spi_data_out_r_39__N_2104[18] (spi_data_out_r_39__N_2104[18]), 
            .\spi_data_out_r_39__N_2249[18] (spi_data_out_r_39__N_2249[18]), 
            .\spi_data_out_r_39__N_2104[17] (spi_data_out_r_39__N_2104[17]), 
            .\spi_data_out_r_39__N_2249[17] (spi_data_out_r_39__N_2249[17]), 
            .\spi_data_out_r_39__N_2104[16] (spi_data_out_r_39__N_2104[16]), 
            .\spi_data_out_r_39__N_2249[16] (spi_data_out_r_39__N_2249[16]), 
            .\spi_data_out_r_39__N_2104[15] (spi_data_out_r_39__N_2104[15]), 
            .\spi_data_out_r_39__N_2249[15] (spi_data_out_r_39__N_2249[15]), 
            .\spi_data_out_r_39__N_2104[14] (spi_data_out_r_39__N_2104[14]), 
            .\spi_data_out_r_39__N_2249[14] (spi_data_out_r_39__N_2249[14]), 
            .\spi_data_out_r_39__N_2104[13] (spi_data_out_r_39__N_2104[13]), 
            .\spi_data_out_r_39__N_2249[13] (spi_data_out_r_39__N_2249[13]), 
            .\spi_data_out_r_39__N_2104[12] (spi_data_out_r_39__N_2104[12]), 
            .\spi_data_out_r_39__N_2249[12] (spi_data_out_r_39__N_2249[12]), 
            .\spi_data_out_r_39__N_2104[11] (spi_data_out_r_39__N_2104[11]), 
            .\spi_data_out_r_39__N_2249[11] (spi_data_out_r_39__N_2249[11]), 
            .\spi_data_out_r_39__N_2104[10] (spi_data_out_r_39__N_2104[10]), 
            .\spi_data_out_r_39__N_2249[10] (spi_data_out_r_39__N_2249[10]), 
            .\spi_data_out_r_39__N_2104[9] (spi_data_out_r_39__N_2104[9]), 
            .\spi_data_out_r_39__N_2249[9] (spi_data_out_r_39__N_2249[9]), 
            .\spi_data_out_r_39__N_2104[8] (spi_data_out_r_39__N_2104[8]), 
            .\spi_data_out_r_39__N_2249[8] (spi_data_out_r_39__N_2249[8]), 
            .\spi_data_out_r_39__N_2104[7] (spi_data_out_r_39__N_2104[7]), 
            .\spi_data_out_r_39__N_2249[7] (spi_data_out_r_39__N_2249[7]), 
            .\spi_data_out_r_39__N_2104[6] (spi_data_out_r_39__N_2104[6]), 
            .\spi_data_out_r_39__N_2249[6] (spi_data_out_r_39__N_2249[6]), 
            .\spi_data_out_r_39__N_2104[5] (spi_data_out_r_39__N_2104[5]), 
            .\spi_data_out_r_39__N_2249[5] (spi_data_out_r_39__N_2249[5]), 
            .\spi_data_out_r_39__N_2104[4] (spi_data_out_r_39__N_2104[4]), 
            .\spi_data_out_r_39__N_2249[4] (spi_data_out_r_39__N_2249[4]), 
            .\spi_data_out_r_39__N_2104[3] (spi_data_out_r_39__N_2104[3]), 
            .\spi_data_out_r_39__N_2249[3] (spi_data_out_r_39__N_2249[3]), 
            .\spi_data_out_r_39__N_2104[2] (spi_data_out_r_39__N_2104[2]), 
            .\spi_data_out_r_39__N_2249[2] (spi_data_out_r_39__N_2249[2]), 
            .\spi_data_out_r_39__N_2104[1] (spi_data_out_r_39__N_2104[1]), 
            .\spi_data_out_r_39__N_2249[1] (spi_data_out_r_39__N_2249[1]), 
            .resetn_c(resetn_c), .GND_net(GND_net), .clk_enable_519(clk_enable_519), 
            .n29079(n29079), .n21446(n21446)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(272[3] 293[2])
    LUT4 m1_lut (.Z(n29757)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    \stepper(DEV_ID=2,UART_ADDRESS_WIDTH=4)  \stepper_ins_2..u_stepper  (.clk_1MHz(clk_1MHz), 
            .clk_1MHz_enable_24(clk_1MHz_enable_24), .n29239(n29239), .mode_adj_134({n29782}), 
            .clk(clk), .clk_enable_271(clk_enable_271), .n29762(n29762), 
            .pin_io_out_29(pin_io_out_29), .\quad_b[2] (quad_b[2]), .pin_io_out_28(pin_io_out_28), 
            .\quad_a[2] (quad_a[2]), .spi_data_out_r_39__N_4496({spi_data_out_r_39__N_4496}), 
            .n47(n47), .digital_output_r(digital_output_r_adj_7976), .clk_enable_190(clk_enable_190), 
            .\spi_data_r[0] (spi_data_r[0]), .n29295(n29295), .spi_data_out_r_39__N_4536(spi_data_out_r_39__N_4536), 
            .n19361(n19361), .resetn_c(resetn_c), .mode(mode_adj_8138), 
            .n29303(n29303), .n22(n22_adj_7754), .GND_net(GND_net), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[1] (spi_data_r[1]), .n1(n1_adj_8169), .n8767(n8767), 
            .n29193(n29193), .reset_r(reset_r_adj_7975), .clk_enable_306(clk_enable_306), 
            .n29070(n29070), .n1_adj_133(n1_adj_8168), .n29117(n29117), 
            .\spi_cmd[2] (spi_cmd[2]), .n29212(n29212), .n13413(n13413), 
            .quad_homing({quad_homing_adj_8284}), .pin_io_out_24(pin_io_out_24), 
            .n29233(n29233), .n12714(n12714)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(364[3] 407[2])
    \stepper(UART_ADDRESS_WIDTH=4)  \stepper_ins_0..u_stepper  (.\spi_cmd[0] (spi_cmd[0]), 
            .n29108(n29108), .\SLO_buf[4] (SLO_buf_adj_8920[4]), .\SLO_buf[14] (SLO_buf_adj_8920[14]), 
            .\spi_data_out_r_39__N_5775[0] (spi_data_out_r_39__N_5775[0]), 
            .\SLO_buf[3] (SLO_buf_adj_8920[3]), .\SLO_buf[9] (SLO_buf_adj_8920[9]), 
            .\spi_data_out_r_39__N_5775[35] (spi_data_out_r_39__N_5775[35]), 
            .\SLO_buf[2] (SLO_buf_adj_8920[2]), .\SLO_buf[8] (SLO_buf_adj_8920[8]), 
            .\spi_data_out_r_39__N_5775[34] (spi_data_out_r_39__N_5775[34]), 
            .\SLO_buf[1] (SLO_buf_adj_8920[1]), .\SLO_buf[7] (SLO_buf_adj_8920[7]), 
            .\spi_data_out_r_39__N_5775[33] (spi_data_out_r_39__N_5775[33]), 
            .n29087(n29087), .\SLO_buf[16] (SLO_buf_adj_8951[16]), .\SLO_buf[26] (SLO_buf_adj_8951[26]), 
            .\spi_data_out_r_39__N_6114[12] (spi_data_out_r_39__N_6114[12]), 
            .\SLO_buf[0] (SLO_buf_adj_8920[0]), .\SLO_buf[6] (SLO_buf_adj_8920[6]), 
            .\spi_data_out_r_39__N_5775[32] (spi_data_out_r_39__N_5775[32]), 
            .\SLO_buf[19] (SLO_buf_adj_8920[19]), .\SLO_buf[29] (SLO_buf_adj_8920[29]), 
            .\spi_data_out_r_39__N_5775[15] (spi_data_out_r_39__N_5775[15]), 
            .\SLO_buf[18] (SLO_buf_adj_8920[18]), .\SLO_buf[28] (SLO_buf_adj_8920[28]), 
            .\spi_data_out_r_39__N_5775[14] (spi_data_out_r_39__N_5775[14]), 
            .\SLO_buf[17] (SLO_buf_adj_8920[17]), .\SLO_buf[27] (SLO_buf_adj_8920[27]), 
            .\spi_data_out_r_39__N_5775[13] (spi_data_out_r_39__N_5775[13]), 
            .\SLO_buf[16]_adj_11 (SLO_buf_adj_8920[16]), .\SLO_buf[26]_adj_12 (SLO_buf_adj_8920[26]), 
            .\spi_data_out_r_39__N_5775[12] (spi_data_out_r_39__N_5775[12]), 
            .\SLO_buf[15] (SLO_buf_adj_8920[15]), .\SLO_buf[25] (SLO_buf_adj_8920[25]), 
            .\spi_data_out_r_39__N_5775[11] (spi_data_out_r_39__N_5775[11]), 
            .\SLO_buf[24] (SLO_buf_adj_8920[24]), .\spi_data_out_r_39__N_5775[10] (spi_data_out_r_39__N_5775[10]), 
            .\SLO_buf[13] (SLO_buf_adj_8920[13]), .\SLO_buf[23] (SLO_buf_adj_8920[23]), 
            .\spi_data_out_r_39__N_5775[9] (spi_data_out_r_39__N_5775[9]), 
            .\SLO_buf[12] (SLO_buf_adj_8920[12]), .\SLO_buf[22] (SLO_buf_adj_8920[22]), 
            .\spi_data_out_r_39__N_5775[8] (spi_data_out_r_39__N_5775[8]), 
            .\SLO_buf[11] (SLO_buf_adj_8920[11]), .\SLO_buf[21] (SLO_buf_adj_8920[21]), 
            .\spi_data_out_r_39__N_5775[7] (spi_data_out_r_39__N_5775[7]), 
            .\SLO_buf[10] (SLO_buf_adj_8920[10]), .\SLO_buf[20] (SLO_buf_adj_8920[20]), 
            .\spi_data_out_r_39__N_5775[6] (spi_data_out_r_39__N_5775[6]), 
            .\spi_data_out_r_39__N_5775[5] (spi_data_out_r_39__N_5775[5]), 
            .\spi_data_out_r_39__N_5775[4] (spi_data_out_r_39__N_5775[4]), 
            .\spi_data_out_r_39__N_5775[3] (spi_data_out_r_39__N_5775[3]), 
            .\spi_data_out_r_39__N_5775[2] (spi_data_out_r_39__N_5775[2]), 
            .pin_io_out_8(pin_io_out_8), .spi_data_out_r_39__N_3818({spi_data_out_r_39__N_3818}), 
            .clk(clk), .\SLO_buf[5] (SLO_buf_adj_8920[5]), .\spi_data_out_r_39__N_5775[1] (spi_data_out_r_39__N_5775[1]), 
            .mode_adj_132({n29780}), .clk_1MHz(clk_1MHz), .n29239(n29239), 
            .pin_io_out_9(pin_io_out_9), .\quad_b[0] (quad_b[0]), .\quad_a[0] (quad_a[0]), 
            .n29201(n29201), .clk_1MHz_enable_55(clk_1MHz_enable_55), .clk_enable_402(clk_enable_402), 
            .n29762(n29762), .n29185(n29185), .\spi_addr[1] (spi_addr[1]), 
            .n29761(n29761), .\spi_addr[2] (spi_addr[2]), .\spi_cmd[2] (spi_cmd[2]), 
            .n13489(n13489), .n29178(n29178), .digital_output_r(digital_output_r), 
            .clk_enable_173(clk_enable_173), .\spi_data_r[0] (spi_data_r[0]), 
            .spi_data_out_r_39__N_3858(spi_data_out_r_39__N_3858), .\SLO_buf[4]_adj_13 (SLO_buf_adj_8951[4]), 
            .\SLO_buf[14]_adj_14 (SLO_buf_adj_8951[14]), .\spi_data_out_r_39__N_6114[0] (spi_data_out_r_39__N_6114[0]), 
            .\SLO_buf[3]_adj_15 (SLO_buf_adj_8951[3]), .\SLO_buf[9]_adj_16 (SLO_buf_adj_8951[9]), 
            .\spi_data_out_r_39__N_6114[35] (spi_data_out_r_39__N_6114[35]), 
            .resetn_c(resetn_c), .n19337(n19337), .\SLO_buf[15]_adj_17 (SLO_buf_adj_8951[15]), 
            .\SLO_buf[25]_adj_18 (SLO_buf_adj_8951[25]), .\spi_data_out_r_39__N_6114[11] (spi_data_out_r_39__N_6114[11]), 
            .\SLO_buf[24]_adj_19 (SLO_buf_adj_8951[24]), .\spi_data_out_r_39__N_6114[10] (spi_data_out_r_39__N_6114[10]), 
            .\SLO_buf[13]_adj_20 (SLO_buf_adj_8951[13]), .\SLO_buf[23]_adj_21 (SLO_buf_adj_8951[23]), 
            .\spi_data_out_r_39__N_6114[9] (spi_data_out_r_39__N_6114[9]), 
            .\SLO_buf[4]_adj_22 (SLO_buf_adj_8889[4]), .\SLO_buf[14]_adj_23 (SLO_buf_adj_8889[14]), 
            .\spi_data_out_r_39__N_5436[0] (spi_data_out_r_39__N_5436[0]), 
            .\SLO_buf[3]_adj_24 (SLO_buf_adj_8889[3]), .\SLO_buf[9]_adj_25 (SLO_buf_adj_8889[9]), 
            .\spi_data_out_r_39__N_5436[35] (spi_data_out_r_39__N_5436[35]), 
            .\SLO_buf[2]_adj_26 (SLO_buf_adj_8951[2]), .\SLO_buf[8]_adj_27 (SLO_buf_adj_8951[8]), 
            .\spi_data_out_r_39__N_6114[34] (spi_data_out_r_39__N_6114[34]), 
            .\SLO_buf[2]_adj_28 (SLO_buf_adj_8889[2]), .\SLO_buf[8]_adj_29 (SLO_buf_adj_8889[8]), 
            .\spi_data_out_r_39__N_5436[34] (spi_data_out_r_39__N_5436[34]), 
            .\SLO_buf[1]_adj_30 (SLO_buf_adj_8889[1]), .\SLO_buf[7]_adj_31 (SLO_buf_adj_8889[7]), 
            .\spi_data_out_r_39__N_5436[33] (spi_data_out_r_39__N_5436[33]), 
            .\SLO_buf[0]_adj_32 (SLO_buf_adj_8889[0]), .\SLO_buf[6]_adj_33 (SLO_buf_adj_8889[6]), 
            .\spi_data_out_r_39__N_5436[32] (spi_data_out_r_39__N_5436[32]), 
            .\SLO_buf[12]_adj_34 (SLO_buf_adj_8951[12]), .\SLO_buf[22]_adj_35 (SLO_buf_adj_8951[22]), 
            .\spi_data_out_r_39__N_6114[8] (spi_data_out_r_39__N_6114[8]), 
            .\SLO_buf[19]_adj_36 (SLO_buf_adj_8889[19]), .\SLO_buf[29]_adj_37 (SLO_buf_adj_8889[29]), 
            .\spi_data_out_r_39__N_5436[15] (spi_data_out_r_39__N_5436[15]), 
            .\SLO_buf[18]_adj_38 (SLO_buf_adj_8889[18]), .\SLO_buf[28]_adj_39 (SLO_buf_adj_8889[28]), 
            .\spi_data_out_r_39__N_5436[14] (spi_data_out_r_39__N_5436[14]), 
            .\SLO_buf[11]_adj_40 (SLO_buf_adj_8951[11]), .\SLO_buf[21]_adj_41 (SLO_buf_adj_8951[21]), 
            .\spi_data_out_r_39__N_6114[7] (spi_data_out_r_39__N_6114[7]), 
            .\SLO_buf[10]_adj_42 (SLO_buf_adj_8951[10]), .\SLO_buf[20]_adj_43 (SLO_buf_adj_8951[20]), 
            .\spi_data_out_r_39__N_6114[6] (spi_data_out_r_39__N_6114[6]), 
            .\SLO_buf[17]_adj_44 (SLO_buf_adj_8889[17]), .\SLO_buf[27]_adj_45 (SLO_buf_adj_8889[27]), 
            .\spi_data_out_r_39__N_5436[13] (spi_data_out_r_39__N_5436[13]), 
            .\SLO_buf[16]_adj_46 (SLO_buf_adj_8889[16]), .\SLO_buf[26]_adj_47 (SLO_buf_adj_8889[26]), 
            .\spi_data_out_r_39__N_5436[12] (spi_data_out_r_39__N_5436[12]), 
            .\SLO_buf[15]_adj_48 (SLO_buf_adj_8889[15]), .\SLO_buf[25]_adj_49 (SLO_buf_adj_8889[25]), 
            .\spi_data_out_r_39__N_5436[11] (spi_data_out_r_39__N_5436[11]), 
            .\SLO_buf[1]_adj_50 (SLO_buf_adj_8951[1]), .\SLO_buf[7]_adj_51 (SLO_buf_adj_8951[7]), 
            .\spi_data_out_r_39__N_6114[33] (spi_data_out_r_39__N_6114[33]), 
            .\SLO_buf[24]_adj_52 (SLO_buf_adj_8889[24]), .\spi_data_out_r_39__N_5436[10] (spi_data_out_r_39__N_5436[10]), 
            .\SLO_buf[13]_adj_53 (SLO_buf_adj_8889[13]), .\SLO_buf[23]_adj_54 (SLO_buf_adj_8889[23]), 
            .\spi_data_out_r_39__N_5436[9] (spi_data_out_r_39__N_5436[9]), 
            .n1(n1_adj_8177), .\SLO_buf[0]_adj_55 (SLO_buf_adj_8951[0]), 
            .\SLO_buf[6]_adj_56 (SLO_buf_adj_8951[6]), .\spi_data_out_r_39__N_6114[32] (spi_data_out_r_39__N_6114[32]), 
            .n29309(n29309), .n8823(n8823), .n29216(n29216), .n29205(n29205), 
            .\spi_addr_r[1] (spi_addr_r[1]), .n29214(n29214), .n29134(n29134), 
            .\SLO_buf[12]_adj_57 (SLO_buf_adj_8889[12]), .\SLO_buf[22]_adj_58 (SLO_buf_adj_8889[22]), 
            .\spi_data_out_r_39__N_5436[8] (spi_data_out_r_39__N_5436[8]), 
            .\SLO_buf[11]_adj_59 (SLO_buf_adj_8889[11]), .\SLO_buf[21]_adj_60 (SLO_buf_adj_8889[21]), 
            .\spi_data_out_r_39__N_5436[7] (spi_data_out_r_39__N_5436[7]), 
            .\SLO_buf[10]_adj_61 (SLO_buf_adj_8889[10]), .\SLO_buf[20]_adj_62 (SLO_buf_adj_8889[20]), 
            .\spi_data_out_r_39__N_5436[6] (spi_data_out_r_39__N_5436[6]), 
            .\spi_data_out_r_39__N_5436[5] (spi_data_out_r_39__N_5436[5]), 
            .\spi_data_out_r_39__N_5436[4] (spi_data_out_r_39__N_5436[4]), 
            .\spi_data_out_r_39__N_5436[3] (spi_data_out_r_39__N_5436[3]), 
            .\spi_data_out_r_39__N_5436[2] (spi_data_out_r_39__N_5436[2]), 
            .\SLO_buf[19]_adj_63 (SLO_buf_adj_8951[19]), .\SLO_buf[29]_adj_64 (SLO_buf_adj_8951[29]), 
            .\spi_data_out_r_39__N_6114[15] (spi_data_out_r_39__N_6114[15]), 
            .n1_adj_65(n1_adj_8176), .\cs_decoded[0] (cs_decoded[0]), .n8824(n8824), 
            .\SLO_buf[5]_adj_66 (SLO_buf_adj_8889[5]), .\spi_data_out_r_39__N_5436[1] (spi_data_out_r_39__N_5436[1]), 
            .\spi_data_out_r_39__N_6114[5] (spi_data_out_r_39__N_6114[5]), 
            .n18550(n18550), .\SLO_buf[18]_adj_67 (SLO_buf_adj_8951[18]), 
            .\spi_data_out_r_39__N_6114[4] (spi_data_out_r_39__N_6114[4]), 
            .GND_net(GND_net), .n29310(n29310), .\SLO_buf[4]_adj_68 (SLO_buf_adj_8858[4]), 
            .\SLO_buf[14]_adj_69 (SLO_buf_adj_8858[14]), .\spi_data_out_r_39__N_5097[0] (spi_data_out_r_39__N_5097[0]), 
            .\SLO_buf[3]_adj_70 (SLO_buf_adj_8858[3]), .\SLO_buf[9]_adj_71 (SLO_buf_adj_8858[9]), 
            .\spi_data_out_r_39__N_5097[35] (spi_data_out_r_39__N_5097[35]), 
            .\SLO_buf[2]_adj_72 (SLO_buf_adj_8858[2]), .\SLO_buf[8]_adj_73 (SLO_buf_adj_8858[8]), 
            .\spi_data_out_r_39__N_5097[34] (spi_data_out_r_39__N_5097[34]), 
            .\SLO_buf[17]_adj_74 (SLO_buf_adj_8951[17]), .\spi_data_out_r_39__N_6114[3] (spi_data_out_r_39__N_6114[3]), 
            .\spi_data_out_r_39__N_6114[2] (spi_data_out_r_39__N_6114[2]), 
            .\SLO_buf[28]_adj_75 (SLO_buf_adj_8951[28]), .\spi_data_out_r_39__N_6114[14] (spi_data_out_r_39__N_6114[14]), 
            .mode(mode_adj_8128), .n31(n31_adj_8085), .n22(n22), .\SLO_buf[1]_adj_76 (SLO_buf_adj_8858[1]), 
            .\SLO_buf[7]_adj_77 (SLO_buf_adj_8858[7]), .\spi_data_out_r_39__N_5097[33] (spi_data_out_r_39__N_5097[33]), 
            .\SLO_buf[0]_adj_78 (SLO_buf_adj_8858[0]), .\SLO_buf[6]_adj_79 (SLO_buf_adj_8858[6]), 
            .\spi_data_out_r_39__N_5097[32] (spi_data_out_r_39__N_5097[32]), 
            .\SLO_buf[5]_adj_80 (SLO_buf_adj_8951[5]), .\spi_data_out_r_39__N_6114[1] (spi_data_out_r_39__N_6114[1]), 
            .\SLO_buf[19]_adj_81 (SLO_buf_adj_8858[19]), .\SLO_buf[29]_adj_82 (SLO_buf_adj_8858[29]), 
            .\spi_data_out_r_39__N_5097[15] (spi_data_out_r_39__N_5097[15]), 
            .\SLO_buf[18]_adj_83 (SLO_buf_adj_8858[18]), .\SLO_buf[28]_adj_84 (SLO_buf_adj_8858[28]), 
            .\spi_data_out_r_39__N_5097[14] (spi_data_out_r_39__N_5097[14]), 
            .\SLO_buf[17]_adj_85 (SLO_buf_adj_8858[17]), .\SLO_buf[27]_adj_86 (SLO_buf_adj_8858[27]), 
            .\spi_data_out_r_39__N_5097[13] (spi_data_out_r_39__N_5097[13]), 
            .\SLO_buf[16]_adj_87 (SLO_buf_adj_8858[16]), .\SLO_buf[26]_adj_88 (SLO_buf_adj_8858[26]), 
            .\spi_data_out_r_39__N_5097[12] (spi_data_out_r_39__N_5097[12]), 
            .\SLO_buf[15]_adj_89 (SLO_buf_adj_8858[15]), .\SLO_buf[25]_adj_90 (SLO_buf_adj_8858[25]), 
            .\spi_data_out_r_39__N_5097[11] (spi_data_out_r_39__N_5097[11]), 
            .\SLO_buf[24]_adj_91 (SLO_buf_adj_8858[24]), .\spi_data_out_r_39__N_5097[10] (spi_data_out_r_39__N_5097[10]), 
            .\SLO_buf[13]_adj_92 (SLO_buf_adj_8858[13]), .\SLO_buf[23]_adj_93 (SLO_buf_adj_8858[23]), 
            .\spi_data_out_r_39__N_5097[9] (spi_data_out_r_39__N_5097[9]), 
            .\SLO_buf[12]_adj_94 (SLO_buf_adj_8858[12]), .\SLO_buf[22]_adj_95 (SLO_buf_adj_8858[22]), 
            .\spi_data_out_r_39__N_5097[8] (spi_data_out_r_39__N_5097[8]), 
            .\SLO_buf[11]_adj_96 (SLO_buf_adj_8858[11]), .\SLO_buf[21]_adj_97 (SLO_buf_adj_8858[21]), 
            .\spi_data_out_r_39__N_5097[7] (spi_data_out_r_39__N_5097[7]), 
            .\SLO_buf[10]_adj_98 (SLO_buf_adj_8858[10]), .\SLO_buf[20]_adj_99 (SLO_buf_adj_8858[20]), 
            .\spi_data_out_r_39__N_5097[6] (spi_data_out_r_39__N_5097[6]), 
            .\spi_cmd_r[1] (spi_cmd_r[1]), .\spi_addr_r[0] (spi_addr_r[0]), 
            .n29287(n29287), .\spi_cmd_r[0] (spi_cmd_r[0]), .n29311(n29311), 
            .n27286(n27286), .\SLO_buf[27]_adj_100 (SLO_buf_adj_8951[27]), 
            .\spi_data_out_r_39__N_6114[13] (spi_data_out_r_39__N_6114[13]), 
            .\spi_data_out_r_39__N_5097[5] (spi_data_out_r_39__N_5097[5]), 
            .\spi_data_out_r_39__N_5097[4] (spi_data_out_r_39__N_5097[4]), 
            .\spi_data_out_r_39__N_5097[3] (spi_data_out_r_39__N_5097[3]), 
            .\spi_data_out_r_39__N_5097[2] (spi_data_out_r_39__N_5097[2]), 
            .\SLO_buf[5]_adj_101 (SLO_buf_adj_8858[5]), .\spi_data_out_r_39__N_5097[1] (spi_data_out_r_39__N_5097[1]), 
            .\SLO_buf[3]_adj_102 (SLO_buf_adj_8796[3]), .\SLO_buf[9]_adj_103 (SLO_buf_adj_8796[9]), 
            .\spi_data_out_r_39__N_4419[35] (spi_data_out_r_39__N_4419[35]), 
            .\SLO_buf[2]_adj_104 (SLO_buf_adj_8796[2]), .\SLO_buf[8]_adj_105 (SLO_buf_adj_8796[8]), 
            .\spi_data_out_r_39__N_4419[34] (spi_data_out_r_39__N_4419[34]), 
            .\SLO_buf[1]_adj_106 (SLO_buf_adj_8796[1]), .\SLO_buf[7]_adj_107 (SLO_buf_adj_8796[7]), 
            .\spi_data_out_r_39__N_4419[33] (spi_data_out_r_39__N_4419[33]), 
            .\SLO_buf[0]_adj_108 (SLO_buf_adj_8796[0]), .\SLO_buf[6]_adj_109 (SLO_buf_adj_8796[6]), 
            .\spi_data_out_r_39__N_4419[32] (spi_data_out_r_39__N_4419[32]), 
            .\SLO_buf[19]_adj_110 (SLO_buf_adj_8796[19]), .\SLO_buf[29]_adj_111 (SLO_buf_adj_8796[29]), 
            .\spi_data_out_r_39__N_4419[15] (spi_data_out_r_39__N_4419[15]), 
            .\SLO_buf[18]_adj_112 (SLO_buf_adj_8796[18]), .\SLO_buf[28]_adj_113 (SLO_buf_adj_8796[28]), 
            .\spi_data_out_r_39__N_4419[14] (spi_data_out_r_39__N_4419[14]), 
            .\SLO_buf[17]_adj_114 (SLO_buf_adj_8796[17]), .\SLO_buf[27]_adj_115 (SLO_buf_adj_8796[27]), 
            .\spi_data_out_r_39__N_4419[13] (spi_data_out_r_39__N_4419[13]), 
            .\SLO_buf[16]_adj_116 (SLO_buf_adj_8796[16]), .\SLO_buf[26]_adj_117 (SLO_buf_adj_8796[26]), 
            .\spi_data_out_r_39__N_4419[12] (spi_data_out_r_39__N_4419[12]), 
            .\SLO_buf[15]_adj_118 (SLO_buf_adj_8796[15]), .\SLO_buf[25]_adj_119 (SLO_buf_adj_8796[25]), 
            .\spi_data_out_r_39__N_4419[11] (spi_data_out_r_39__N_4419[11]), 
            .\SLO_buf[14]_adj_120 (SLO_buf_adj_8796[14]), .\SLO_buf[24]_adj_121 (SLO_buf_adj_8796[24]), 
            .\spi_data_out_r_39__N_4419[10] (spi_data_out_r_39__N_4419[10]), 
            .\SLO_buf[13]_adj_122 (SLO_buf_adj_8796[13]), .\SLO_buf[23]_adj_123 (SLO_buf_adj_8796[23]), 
            .\spi_data_out_r_39__N_4419[9] (spi_data_out_r_39__N_4419[9]), 
            .\SLO_buf[12]_adj_124 (SLO_buf_adj_8796[12]), .\SLO_buf[22]_adj_125 (SLO_buf_adj_8796[22]), 
            .\spi_data_out_r_39__N_4419[8] (spi_data_out_r_39__N_4419[8]), 
            .\SLO_buf[11]_adj_126 (SLO_buf_adj_8796[11]), .\SLO_buf[21]_adj_127 (SLO_buf_adj_8796[21]), 
            .\spi_data_out_r_39__N_4419[7] (spi_data_out_r_39__N_4419[7]), 
            .\SLO_buf[10]_adj_128 (SLO_buf_adj_8796[10]), .\SLO_buf[20]_adj_129 (SLO_buf_adj_8796[20]), 
            .\spi_data_out_r_39__N_4419[6] (spi_data_out_r_39__N_4419[6]), 
            .\spi_data_out_r_39__N_4419[5] (spi_data_out_r_39__N_4419[5]), 
            .\spi_data_out_r_39__N_4419[4] (spi_data_out_r_39__N_4419[4]), 
            .\spi_data_out_r_39__N_4419[3] (spi_data_out_r_39__N_4419[3]), 
            .\spi_data_out_r_39__N_4419[2] (spi_data_out_r_39__N_4419[2]), 
            .\SLO_buf[5]_adj_130 (SLO_buf_adj_8796[5]), .\spi_data_out_r_39__N_4419[1] (spi_data_out_r_39__N_4419[1]), 
            .\SLO_buf[4]_adj_131 (SLO_buf_adj_8796[4]), .\spi_data_out_r_39__N_4419[0] (spi_data_out_r_39__N_4419[0]), 
            .\spi_data_r[1] (spi_data_r[1]), .\spi_data_r[2] (spi_data_r[2]), 
            .reset_r(reset_r), .clk_enable_506(clk_enable_506), .n29106(n29106), 
            .n29117(n29117), .n29076(n29076), .n29115(n29115), .spi_data_out_r_39__N_4490(spi_data_out_r_39__N_4490), 
            .n29093(n29093), .n29094(n29094), .\spi_addr[0] (spi_addr[0]), 
            .n29126(n29126), .clear_intrpt_N_2710(clear_intrpt_N_2710), 
            .\spi_cmd[1] (spi_cmd[1]), .n29141(n29141), .n26933(n26933), 
            .n29212(n29212), .n47(n47), .clear_intrpt_N_2639(clear_intrpt_N_2639), 
            .spi_data_out_r_39__N_5507(spi_data_out_r_39__N_5507), .n29091(n29091), 
            .n29098(n29098), .n29099(n29099)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(364[3] 407[2])
    \stepper(DEV_ID=4,UART_ADDRESS_WIDTH=4)  \stepper_ins_4..u_stepper  (.GND_net(GND_net), 
            .clk_1MHz(clk_1MHz), .clk_1MHz_enable_66(clk_1MHz_enable_66), 
            .n29239(n29239), .\SLO_buf[0] (SLO_buf_adj_8889[0]), .pin_io_out_48(pin_io_out_48), 
            .spi_data_out_r_39__N_5174({spi_data_out_r_39__N_5174}), .clk(clk), 
            .\spi_data_out_r_39__N_5436[0] (spi_data_out_r_39__N_5436[0]), 
            .mode_adj_10({n29784}), .clk_enable_359(clk_enable_359), .n29762(n29762), 
            .n29091(n29091), .\SLO_buf[13] (SLO_buf_adj_8889[13]), .\SLO_buf[12] (SLO_buf_adj_8889[12]), 
            .\SLO_buf[11] (SLO_buf_adj_8889[11]), .\SLO_buf[10] (SLO_buf_adj_8889[10]), 
            .\spi_data_out_r_39__N_5436[35] (spi_data_out_r_39__N_5436[35]), 
            .\spi_data_out_r_39__N_5436[34] (spi_data_out_r_39__N_5436[34]), 
            .\spi_data_out_r_39__N_5436[33] (spi_data_out_r_39__N_5436[33]), 
            .\spi_data_out_r_39__N_5436[32] (spi_data_out_r_39__N_5436[32]), 
            .\spi_data_out_r_39__N_5436[15] (spi_data_out_r_39__N_5436[15]), 
            .\spi_data_out_r_39__N_5436[14] (spi_data_out_r_39__N_5436[14]), 
            .\spi_data_out_r_39__N_5436[13] (spi_data_out_r_39__N_5436[13]), 
            .\spi_data_out_r_39__N_5436[12] (spi_data_out_r_39__N_5436[12]), 
            .\spi_data_out_r_39__N_5436[11] (spi_data_out_r_39__N_5436[11]), 
            .\spi_data_out_r_39__N_5436[10] (spi_data_out_r_39__N_5436[10]), 
            .\spi_data_out_r_39__N_5436[9] (spi_data_out_r_39__N_5436[9]), 
            .\spi_data_out_r_39__N_5436[8] (spi_data_out_r_39__N_5436[8]), 
            .\spi_data_out_r_39__N_5436[7] (spi_data_out_r_39__N_5436[7]), 
            .\spi_data_out_r_39__N_5436[6] (spi_data_out_r_39__N_5436[6]), 
            .\spi_data_out_r_39__N_5436[5] (spi_data_out_r_39__N_5436[5]), 
            .\spi_data_out_r_39__N_5436[4] (spi_data_out_r_39__N_5436[4]), 
            .\spi_data_out_r_39__N_5436[3] (spi_data_out_r_39__N_5436[3]), 
            .\spi_data_out_r_39__N_5436[2] (spi_data_out_r_39__N_5436[2]), 
            .\spi_data_out_r_39__N_5436[1] (spi_data_out_r_39__N_5436[1]), 
            .\SLO_buf[29] (SLO_buf_adj_8889[29]), .\SLO_buf[28] (SLO_buf_adj_8889[28]), 
            .\SLO_buf[27] (SLO_buf_adj_8889[27]), .\SLO_buf[26] (SLO_buf_adj_8889[26]), 
            .\SLO_buf[25] (SLO_buf_adj_8889[25]), .\SLO_buf[24] (SLO_buf_adj_8889[24]), 
            .\SLO_buf[23] (SLO_buf_adj_8889[23]), .\SLO_buf[22] (SLO_buf_adj_8889[22]), 
            .\SLO_buf[21] (SLO_buf_adj_8889[21]), .\SLO_buf[20] (SLO_buf_adj_8889[20]), 
            .\SLO_buf[19] (SLO_buf_adj_8889[19]), .\SLO_buf[18] (SLO_buf_adj_8889[18]), 
            .\SLO_buf[17] (SLO_buf_adj_8889[17]), .\SLO_buf[16] (SLO_buf_adj_8889[16]), 
            .\SLO_buf[15] (SLO_buf_adj_8889[15]), .\SLO_buf[14] (SLO_buf_adj_8889[14]), 
            .\SLO_buf[9] (SLO_buf_adj_8889[9]), .\SLO_buf[8] (SLO_buf_adj_8889[8]), 
            .\SLO_buf[7] (SLO_buf_adj_8889[7]), .\SLO_buf[6] (SLO_buf_adj_8889[6]), 
            .\SLO_buf[5] (SLO_buf_adj_8889[5]), .\SLO_buf[4] (SLO_buf_adj_8889[4]), 
            .\SLO_buf[3] (SLO_buf_adj_8889[3]), .\SLO_buf[2] (SLO_buf_adj_8889[2]), 
            .\SLO_buf[1] (SLO_buf_adj_8889[1]), .spi_data_out_r_39__N_5214(spi_data_out_r_39__N_5214), 
            .spi_data_out_r_39__N_5507(spi_data_out_r_39__N_5507), .digital_output_r(digital_output_r_adj_8018), 
            .clk_enable_206(clk_enable_206), .\spi_data_r[0] (spi_data_r[0]), 
            .n29207(n29207), .n29189(n29189), .n5(n5), .C_5_c_c(C_5_c_c), 
            .n26965(n26965), .n19381(n19381), .resetn_c(resetn_c), .n29204(n29204), 
            .OW_ID_N_5482(OW_ID_N_5482), .n29285(n29285), .mode(mode_adj_8140), 
            .n27477(n27477), .n25411(n25411), .pin_io_out_49(pin_io_out_49), 
            .\quad_b[4] (quad_b[4]), .\quad_a[4] (quad_a[4]), .n1(n1_adj_8162), 
            .n1_adj_9(n1_adj_8161), .\spi_data_r[1] (spi_data_r[1]), .\spi_data_r[2] (spi_data_r[2]), 
            .pin_io_out_44(pin_io_out_44), .n29224(n29224), .quad_homing({quad_homing_adj_8402}), 
            .n26938(n26938), .reset_r(reset_r_adj_8017), .clk_enable_526(clk_enable_526), 
            .n29077(n29077)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(364[3] 407[2])
    VLO i1 (.Z(GND_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    \rs232(DEV_ID=4,UART_ADDRESS_WIDTH=4)  u_rs232 (.\spi_addr_r[0] (spi_addr_r[0]), 
            .\spi_cmd_r[1] (spi_cmd_r[1]), .n29255(n29255), .n29256(n29256), 
            .n65(n65_adj_8152), .n29083(n29083), .clk(clk), .clk_enable_200(clk_enable_200), 
            .n29239(n29239), .\spi_data_r[0] (spi_data_r[0]), .C_3_c_2(C_3_c_2), 
            .n29282(n29282), .C_4_c_3(C_4_c_3), .n29189(n29189)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(552[3] 572[2])
    \stepper(DEV_ID=1,UART_ADDRESS_WIDTH=4)  \stepper_ins_1..u_stepper  (.mode({n29781}), 
            .clk(clk), .clk_enable_30(clk_enable_30), .n29239(n29239), 
            .\spi_data_r[2] (spi_data_r[2]), .\spi_data_r[1] (spi_data_r[1]), 
            .digital_output_r(digital_output_r_adj_7970), .clk_enable_20(clk_enable_20), 
            .\spi_data_r[0] (spi_data_r[0]), .spi_data_out_r_39__N_4157({spi_data_out_r_39__N_4157}), 
            .n29094(n29094), .\SLO_buf[13] (SLO_buf_adj_8796[13]), .\SLO_buf[12] (SLO_buf_adj_8796[12]), 
            .\SLO_buf[11] (SLO_buf_adj_8796[11]), .\SLO_buf[10] (SLO_buf_adj_8796[10]), 
            .\spi_data_out_r_39__N_4419[35] (spi_data_out_r_39__N_4419[35]), 
            .\spi_data_out_r_39__N_4419[34] (spi_data_out_r_39__N_4419[34]), 
            .\spi_data_out_r_39__N_4419[33] (spi_data_out_r_39__N_4419[33]), 
            .\spi_data_out_r_39__N_4419[32] (spi_data_out_r_39__N_4419[32]), 
            .\spi_data_out_r_39__N_4419[15] (spi_data_out_r_39__N_4419[15]), 
            .\spi_data_out_r_39__N_4419[14] (spi_data_out_r_39__N_4419[14]), 
            .\spi_data_out_r_39__N_4419[13] (spi_data_out_r_39__N_4419[13]), 
            .\spi_data_out_r_39__N_4419[12] (spi_data_out_r_39__N_4419[12]), 
            .\spi_data_out_r_39__N_4419[11] (spi_data_out_r_39__N_4419[11]), 
            .\spi_data_out_r_39__N_4419[10] (spi_data_out_r_39__N_4419[10]), 
            .\spi_data_out_r_39__N_4419[9] (spi_data_out_r_39__N_4419[9]), 
            .\spi_data_out_r_39__N_4419[8] (spi_data_out_r_39__N_4419[8]), 
            .\spi_data_out_r_39__N_4419[7] (spi_data_out_r_39__N_4419[7]), 
            .\spi_data_out_r_39__N_4419[6] (spi_data_out_r_39__N_4419[6]), 
            .\spi_data_out_r_39__N_4419[5] (spi_data_out_r_39__N_4419[5]), 
            .\spi_data_out_r_39__N_4419[4] (spi_data_out_r_39__N_4419[4]), 
            .\spi_data_out_r_39__N_4419[3] (spi_data_out_r_39__N_4419[3]), 
            .\spi_data_out_r_39__N_4419[2] (spi_data_out_r_39__N_4419[2]), 
            .\spi_data_out_r_39__N_4419[1] (spi_data_out_r_39__N_4419[1]), 
            .pin_io_out_19(pin_io_out_19), .\quad_b[1] (quad_b[1]), .pin_io_out_18(pin_io_out_18), 
            .\quad_a[1] (quad_a[1]), .GND_net(GND_net), .clk_1MHz(clk_1MHz), 
            .clk_1MHz_enable_91(clk_1MHz_enable_91), .\SLO_buf[0] (SLO_buf_adj_8796[0]), 
            .\spi_data_out_r_39__N_4419[0] (spi_data_out_r_39__N_4419[0]), 
            .spi_data_out_r_39__N_4197(spi_data_out_r_39__N_4197), .spi_data_out_r_39__N_4490(spi_data_out_r_39__N_4490), 
            .n29762(n29762), .\SLO_buf[29] (SLO_buf_adj_8796[29]), .\SLO_buf[28] (SLO_buf_adj_8796[28]), 
            .\SLO_buf[27] (SLO_buf_adj_8796[27]), .\SLO_buf[26] (SLO_buf_adj_8796[26]), 
            .\SLO_buf[25] (SLO_buf_adj_8796[25]), .\SLO_buf[24] (SLO_buf_adj_8796[24]), 
            .\SLO_buf[23] (SLO_buf_adj_8796[23]), .\SLO_buf[22] (SLO_buf_adj_8796[22]), 
            .\SLO_buf[21] (SLO_buf_adj_8796[21]), .\SLO_buf[20] (SLO_buf_adj_8796[20]), 
            .\SLO_buf[19] (SLO_buf_adj_8796[19]), .\SLO_buf[18] (SLO_buf_adj_8796[18]), 
            .\SLO_buf[17] (SLO_buf_adj_8796[17]), .\SLO_buf[16] (SLO_buf_adj_8796[16]), 
            .\SLO_buf[15] (SLO_buf_adj_8796[15]), .\SLO_buf[14] (SLO_buf_adj_8796[14]), 
            .\SLO_buf[9] (SLO_buf_adj_8796[9]), .\SLO_buf[8] (SLO_buf_adj_8796[8]), 
            .\SLO_buf[7] (SLO_buf_adj_8796[7]), .\SLO_buf[6] (SLO_buf_adj_8796[6]), 
            .\SLO_buf[5] (SLO_buf_adj_8796[5]), .\SLO_buf[4] (SLO_buf_adj_8796[4]), 
            .\SLO_buf[3] (SLO_buf_adj_8796[3]), .\SLO_buf[2] (SLO_buf_adj_8796[2]), 
            .\SLO_buf[1] (SLO_buf_adj_8796[1]), .n19351(n19351), .resetn_c(resetn_c), 
            .n29217(n29217), .n29315(n29315), .\cs_decoded[2] (cs_decoded[2]), 
            .n29306(n29306), .n8796(n8796), .OW_ID_N_4464(OW_ID_N_4464), 
            .C_5_c_c(C_5_c_c), .OW_ID_N_4462(OW_ID_N_4462), .reset_r(reset_r_adj_7969), 
            .clk_enable_307(clk_enable_307), .n29097(n29097), .n1(n1_adj_8173), 
            .n1_adj_8(n1_adj_8172)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(364[3] 407[2])
    \stepper(DEV_ID=5,UART_ADDRESS_WIDTH=4)  \stepper_ins_5..u_stepper  (.\SLO_buf[29] (SLO_buf_adj_8920[29]), 
            .\SLO_buf[28] (SLO_buf_adj_8920[28]), .\SLO_buf[27] (SLO_buf_adj_8920[27]), 
            .\SLO_buf[26] (SLO_buf_adj_8920[26]), .\SLO_buf[25] (SLO_buf_adj_8920[25]), 
            .\SLO_buf[24] (SLO_buf_adj_8920[24]), .\SLO_buf[23] (SLO_buf_adj_8920[23]), 
            .\SLO_buf[22] (SLO_buf_adj_8920[22]), .\SLO_buf[21] (SLO_buf_adj_8920[21]), 
            .\SLO_buf[20] (SLO_buf_adj_8920[20]), .\SLO_buf[19] (SLO_buf_adj_8920[19]), 
            .\SLO_buf[18] (SLO_buf_adj_8920[18]), .\SLO_buf[17] (SLO_buf_adj_8920[17]), 
            .\SLO_buf[16] (SLO_buf_adj_8920[16]), .\SLO_buf[15] (SLO_buf_adj_8920[15]), 
            .\SLO_buf[14] (SLO_buf_adj_8920[14]), .\SLO_buf[13] (SLO_buf_adj_8920[13]), 
            .\SLO_buf[12] (SLO_buf_adj_8920[12]), .\SLO_buf[11] (SLO_buf_adj_8920[11]), 
            .\SLO_buf[10] (SLO_buf_adj_8920[10]), .\SLO_buf[9] (SLO_buf_adj_8920[9]), 
            .\SLO_buf[8] (SLO_buf_adj_8920[8]), .\SLO_buf[7] (SLO_buf_adj_8920[7]), 
            .\SLO_buf[6] (SLO_buf_adj_8920[6]), .\SLO_buf[5] (SLO_buf_adj_8920[5]), 
            .\SLO_buf[4] (SLO_buf_adj_8920[4]), .\SLO_buf[3] (SLO_buf_adj_8920[3]), 
            .\SLO_buf[2] (SLO_buf_adj_8920[2]), .\SLO_buf[1] (SLO_buf_adj_8920[1]), 
            .clk_1MHz(clk_1MHz), .clk_1MHz_enable_40(clk_1MHz_enable_40), 
            .n29239(n29239), .\SLO_buf[0] (SLO_buf_adj_8920[0]), .pin_io_out_58(pin_io_out_58), 
            .spi_data_out_r_39__N_5513({spi_data_out_r_39__N_5513}), .clk(clk), 
            .\spi_data_out_r_39__N_5775[0] (spi_data_out_r_39__N_5775[0]), 
            .mode_adj_7({n29785}), .clk_enable_400(clk_enable_400), .n29762(n29762), 
            .n19391(n19391), .spi_data_out_r_39__N_5553(spi_data_out_r_39__N_5553), 
            .n29108(n29108), .digital_output_r(digital_output_r_adj_8054), 
            .clk_enable_199(clk_enable_199), .\spi_data_r[0] (spi_data_r[0]), 
            .resetn_c(resetn_c), .n29301(n29301), .n29299(n29299), .\cs_decoded[10] (cs_decoded[10]), 
            .n8680(n8680), .n29210(n29210), .n1(n1_adj_8158), .n1_adj_6(n1_adj_8157), 
            .reset_r(reset_r_adj_8053), .clk_enable_342(clk_enable_342), 
            .n29075(n29075), .n29305(n29305), .\spi_data_out_r_39__N_5775[1] (spi_data_out_r_39__N_5775[1]), 
            .\spi_data_out_r_39__N_5775[2] (spi_data_out_r_39__N_5775[2]), 
            .\spi_data_out_r_39__N_5775[3] (spi_data_out_r_39__N_5775[3]), 
            .\spi_data_out_r_39__N_5775[4] (spi_data_out_r_39__N_5775[4]), 
            .\spi_data_out_r_39__N_5775[5] (spi_data_out_r_39__N_5775[5]), 
            .\spi_data_out_r_39__N_5775[6] (spi_data_out_r_39__N_5775[6]), 
            .\spi_data_out_r_39__N_5775[7] (spi_data_out_r_39__N_5775[7]), 
            .\spi_data_out_r_39__N_5775[8] (spi_data_out_r_39__N_5775[8]), 
            .\spi_data_out_r_39__N_5775[9] (spi_data_out_r_39__N_5775[9]), 
            .\spi_data_out_r_39__N_5775[10] (spi_data_out_r_39__N_5775[10]), 
            .\spi_data_out_r_39__N_5775[11] (spi_data_out_r_39__N_5775[11]), 
            .\spi_data_out_r_39__N_5775[12] (spi_data_out_r_39__N_5775[12]), 
            .\spi_data_out_r_39__N_5775[13] (spi_data_out_r_39__N_5775[13]), 
            .\spi_data_out_r_39__N_5775[14] (spi_data_out_r_39__N_5775[14]), 
            .\spi_data_out_r_39__N_5775[15] (spi_data_out_r_39__N_5775[15]), 
            .\spi_data_out_r_39__N_5775[32] (spi_data_out_r_39__N_5775[32]), 
            .\spi_data_out_r_39__N_5775[33] (spi_data_out_r_39__N_5775[33]), 
            .\spi_data_out_r_39__N_5775[34] (spi_data_out_r_39__N_5775[34]), 
            .\spi_data_out_r_39__N_5775[35] (spi_data_out_r_39__N_5775[35]), 
            .pin_io_out_59(pin_io_out_59), .\quad_b[5] (quad_b[5]), .\quad_a[5] (quad_a[5]), 
            .\spi_data_r[1] (spi_data_r[1]), .\spi_data_r[2] (spi_data_r[2]), 
            .mode(mode_adj_8149), .n6(n6_adj_8121), .n29115(n29115), .n18550(n18550), 
            .\spi_addr[1] (spi_addr[1]), .\spi_cmd[0] (spi_cmd[0]), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(364[3] 407[2])
    \uart_controller(DEV_ID=10,UART_ADDRESS_WIDTH=4)  u_uart_controller (.C_1_c_0(C_1_c_0), 
            .clk(clk), .clk_enable_509(clk_enable_509), .n29239(n29239), 
            .\spi_data_r[0] (spi_data_r[0]), .C_2_c_1(C_2_c_1), .\spi_data_r[1] (spi_data_r[1]), 
            .C_3_c_2(C_3_c_2), .\spi_data_r[2] (spi_data_r[2]), .C_4_c_3(C_4_c_3), 
            .\spi_data_r[3] (spi_data_r[3])) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(252[3] 263[2])
    \piezo(DEV_ID=5,UART_ADDRESS_WIDTH=4)  \piezo_ins_5..u_piezo  (.mode(mode_adj_8149), 
            .clk(clk), .clk_enable_174(clk_enable_174), .n29239(n29239), 
            .\spi_data_r[0] (spi_data_r[0]), .mode_adj_5({n29785}), .digital_output_r(digital_output_r_adj_8054), 
            .n26523(n26523), .n29199(n29199), .mode_adj_3(mode_adj_8141), 
            .n6(n6_adj_8121), .mode_adj_4(mode_adj_8133), .n27186(n27186), 
            .C_3_c_2(C_3_c_2), .C_4_c_3(C_4_c_3), .n29313(n29313), .C_2_c_1(C_2_c_1), 
            .C_1_c_0(C_1_c_0), .n29191(n29191), .\cs_decoded[11] (cs_decoded[11]), 
            .n2(n2_adj_8159), .n8850(n8850), .C_5_c_c(C_5_c_c), .n26579(n26579), 
            .n8840(n8840)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(632[3] 661[2])
    GSR GSR_INST (.GSR(resetn_c));
    \stepper(DEV_ID=3,UART_ADDRESS_WIDTH=4)  \stepper_ins_3..u_stepper  (.mode_adj_2({n29783}), 
            .pin_io_out_38(pin_io_out_38), .\quad_a[3] (quad_a[3]), .clk_1MHz(clk_1MHz), 
            .n29239(n29239), .clk_1MHz_enable_182(clk_1MHz_enable_182), 
            .n29203(n29203), .\SLO_buf[0] (SLO_buf_adj_8858[0]), .spi_data_out_r_39__N_4835({spi_data_out_r_39__N_4835}), 
            .clk(clk), .\spi_data_out_r_39__N_5097[0] (spi_data_out_r_39__N_5097[0]), 
            .clk_enable_86(clk_enable_86), .n29762(n29762), .\spi_data_r[2] (spi_data_r[2]), 
            .\spi_data_r[1] (spi_data_r[1]), .n29093(n29093), .\SLO_buf[13] (SLO_buf_adj_8858[13]), 
            .\SLO_buf[12] (SLO_buf_adj_8858[12]), .\SLO_buf[11] (SLO_buf_adj_8858[11]), 
            .\SLO_buf[10] (SLO_buf_adj_8858[10]), .\spi_data_out_r_39__N_5097[35] (spi_data_out_r_39__N_5097[35]), 
            .\spi_data_out_r_39__N_5097[34] (spi_data_out_r_39__N_5097[34]), 
            .\spi_data_out_r_39__N_5097[33] (spi_data_out_r_39__N_5097[33]), 
            .\spi_data_out_r_39__N_5097[32] (spi_data_out_r_39__N_5097[32]), 
            .\spi_data_out_r_39__N_5097[15] (spi_data_out_r_39__N_5097[15]), 
            .\spi_data_out_r_39__N_5097[14] (spi_data_out_r_39__N_5097[14]), 
            .\spi_data_out_r_39__N_5097[13] (spi_data_out_r_39__N_5097[13]), 
            .\spi_data_out_r_39__N_5097[12] (spi_data_out_r_39__N_5097[12]), 
            .\spi_data_out_r_39__N_5097[11] (spi_data_out_r_39__N_5097[11]), 
            .\spi_data_out_r_39__N_5097[10] (spi_data_out_r_39__N_5097[10]), 
            .\spi_data_out_r_39__N_5097[9] (spi_data_out_r_39__N_5097[9]), 
            .\spi_data_out_r_39__N_5097[8] (spi_data_out_r_39__N_5097[8]), 
            .\spi_data_out_r_39__N_5097[7] (spi_data_out_r_39__N_5097[7]), 
            .\spi_data_out_r_39__N_5097[6] (spi_data_out_r_39__N_5097[6]), 
            .\spi_data_out_r_39__N_5097[5] (spi_data_out_r_39__N_5097[5]), 
            .\spi_data_out_r_39__N_5097[4] (spi_data_out_r_39__N_5097[4]), 
            .\spi_data_out_r_39__N_5097[3] (spi_data_out_r_39__N_5097[3]), 
            .\spi_data_out_r_39__N_5097[2] (spi_data_out_r_39__N_5097[2]), 
            .\spi_data_out_r_39__N_5097[1] (spi_data_out_r_39__N_5097[1]), 
            .n29317(n29317), .\SLO_buf[29] (SLO_buf_adj_8858[29]), .\SLO_buf[28] (SLO_buf_adj_8858[28]), 
            .\SLO_buf[27] (SLO_buf_adj_8858[27]), .\SLO_buf[26] (SLO_buf_adj_8858[26]), 
            .\SLO_buf[25] (SLO_buf_adj_8858[25]), .\SLO_buf[24] (SLO_buf_adj_8858[24]), 
            .\SLO_buf[23] (SLO_buf_adj_8858[23]), .\SLO_buf[22] (SLO_buf_adj_8858[22]), 
            .\SLO_buf[21] (SLO_buf_adj_8858[21]), .\SLO_buf[20] (SLO_buf_adj_8858[20]), 
            .\SLO_buf[19] (SLO_buf_adj_8858[19]), .\SLO_buf[18] (SLO_buf_adj_8858[18]), 
            .\SLO_buf[17] (SLO_buf_adj_8858[17]), .\SLO_buf[16] (SLO_buf_adj_8858[16]), 
            .\SLO_buf[15] (SLO_buf_adj_8858[15]), .\SLO_buf[14] (SLO_buf_adj_8858[14]), 
            .\SLO_buf[9] (SLO_buf_adj_8858[9]), .\SLO_buf[8] (SLO_buf_adj_8858[8]), 
            .\SLO_buf[7] (SLO_buf_adj_8858[7]), .\SLO_buf[6] (SLO_buf_adj_8858[6]), 
            .\SLO_buf[5] (SLO_buf_adj_8858[5]), .\SLO_buf[4] (SLO_buf_adj_8858[4]), 
            .\SLO_buf[3] (SLO_buf_adj_8858[3]), .\SLO_buf[2] (SLO_buf_adj_8858[2]), 
            .\SLO_buf[1] (SLO_buf_adj_8858[1]), .digital_output_r(digital_output_r_adj_7982), 
            .clk_enable_164(clk_enable_164), .\spi_data_r[0] (spi_data_r[0]), 
            .spi_data_out_r_39__N_4875(spi_data_out_r_39__N_4875), .n19371(n19371), 
            .resetn_c(resetn_c), .GND_net(GND_net), .NSL(NSL), .mode(mode_adj_8139), 
            .n29300(n29300), .n29149(n29149), .pin_io_out_39(pin_io_out_39), 
            .\quad_b[3] (quad_b[3]), .reset_r(reset_r_adj_7981), .clk_enable_340(clk_enable_340), 
            .n29110(n29110), .n1(n1_adj_8165), .mode_adj_1(mode_adj_8143), 
            .n8716(n8716), .n29115(n29115), .\spi_cmd[2] (spi_cmd[2]), 
            .n13413(n13413)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/mcm_top.v(364[3] 407[2])
    
endmodule
//
// Verilog Description of module \io(DEV_ID=3,UART_ADDRESS_WIDTH=4) 
//

module \io(DEV_ID=3,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_201, 
            n29239, \spi_data_r[0] ) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_201;
    input n29239;
    input \spi_data_r[0] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    FD1P3IX mode_90 (.D(\spi_data_r[0] ), .SP(clk_enable_201), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=464, LSE_RLINE=496 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(80[8] 88[4])
    defparam mode_90.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \shutter(DEV_ID=3,UART_ADDRESS_WIDTH=4) 
//

module \shutter(DEV_ID=3,UART_ADDRESS_WIDTH=4)  (\mode[1] , \mode[2] , n29225, 
            \quad_homing[1] , n27632, n26969, n13052, pin_io_out_34, 
            \pin_intrpt[11] , pin_io_out_32, \pin_intrpt[9] , reset_r, 
            n1, \cs_decoded[6] , n2, pin_io_out_33, \pin_intrpt[10] , 
            mode, clk, clk_enable_171, n29239, \spi_data_r[0] ) /* synthesis syn_module_defined=1 */ ;
    input \mode[1] ;
    input \mode[2] ;
    output n29225;
    input \quad_homing[1] ;
    input n27632;
    output n26969;
    output n13052;
    input pin_io_out_34;
    output \pin_intrpt[11] ;
    input pin_io_out_32;
    output \pin_intrpt[9] ;
    input reset_r;
    output n1;
    input \cs_decoded[6] ;
    output n2;
    input pin_io_out_33;
    output \pin_intrpt[10] ;
    output mode;
    input clk;
    input clk_enable_171;
    input n29239;
    input \spi_data_r[0] ;
    
    wire \pin_intrpt[11]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[11] */ ;   // c:/s_links/sources/mcm_top.v(102[46:56])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    LUT4 i22745_2_lut_rep_497 (.A(\mode[1] ), .B(\mode[2] ), .Z(n29225)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i22745_2_lut_rep_497.init = 16'h1111;
    LUT4 i2_3_lut_4_lut (.A(\mode[1] ), .B(\mode[2] ), .C(\quad_homing[1] ), 
         .D(n27632), .Z(n26969)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;
    defparam i2_3_lut_4_lut.init = 16'hf1ff;
    LUT4 i3_3_lut_4_lut (.A(\mode[1] ), .B(\mode[2] ), .C(\quad_homing[1] ), 
         .D(n27632), .Z(n13052)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i3_3_lut_4_lut.init = 16'h0e00;
    LUT4 i4192_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(pin_io_out_34), 
         .Z(\pin_intrpt[11] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i4192_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_4108_i1_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(pin_io_out_32), 
         .Z(\pin_intrpt[9] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4108_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_3953_i1_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(reset_r), 
         .Z(n1)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_3953_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_3940_i2_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(\cs_decoded[6] ), 
         .Z(n2)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_3940_i2_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_4107_i1_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(pin_io_out_33), 
         .Z(\pin_intrpt[10] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4107_i1_2_lut_3_lut.init = 16'he0e0;
    FD1P3IX mode_160 (.D(\spi_data_r[0] ), .SP(clk_enable_171), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=508, LSE_RLINE=540 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(81[8] 89[4])
    defparam mode_160.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \shutter(DEV_ID=2,UART_ADDRESS_WIDTH=4) 
//

module \shutter(DEV_ID=2,UART_ADDRESS_WIDTH=4)  (\mode[1] , \mode[2] , n29233, 
            pin_io_out_22, \pin_intrpt[6] , reset_r, n1, \cs_decoded[4] , 
            n2, pin_io_out_24, \mode[2]_derived_32 , pin_io_out_23, 
            \pin_intrpt[7] , mode, clk, clk_enable_176, n29239, \spi_data_r[0] , 
            n29194, n29193, n29303, n27480) /* synthesis syn_module_defined=1 */ ;
    input \mode[1] ;
    input \mode[2] ;
    output n29233;
    input pin_io_out_22;
    output \pin_intrpt[6] ;
    input reset_r;
    output n1;
    input \cs_decoded[4] ;
    output n2;
    input pin_io_out_24;
    output \mode[2]_derived_32 ;
    input pin_io_out_23;
    output \pin_intrpt[7] ;
    output mode;
    input clk;
    input clk_enable_176;
    input n29239;
    input \spi_data_r[0] ;
    input n29194;
    input n29193;
    input n29303;
    output n27480;
    
    wire \mode[2]_derived_32  /* synthesis is_clock=1, SET_AS_NETWORK=\stepper_ins[2].u_stepper/mode[2]_derived_32 */ ;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    LUT4 i22733_2_lut_rep_505 (.A(\mode[1] ), .B(\mode[2] ), .Z(n29233)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i22733_2_lut_rep_505.init = 16'h1111;
    LUT4 Select_4110_i1_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(pin_io_out_22), 
         .Z(\pin_intrpt[6] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4110_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_3982_i1_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(reset_r), 
         .Z(n1)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_3982_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_3969_i2_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(\cs_decoded[4] ), 
         .Z(n2)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_3969_i2_2_lut_3_lut.init = 16'he0e0;
    LUT4 i22409_2_lut_rep_444_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(pin_io_out_24), 
         .Z(\mode[2]_derived_32 )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i22409_2_lut_rep_444_3_lut.init = 16'he0e0;
    LUT4 Select_4109_i1_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(pin_io_out_23), 
         .Z(\pin_intrpt[7] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4109_i1_2_lut_3_lut.init = 16'he0e0;
    FD1P3IX mode_160 (.D(\spi_data_r[0] ), .SP(clk_enable_176), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=508, LSE_RLINE=540 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(81[8] 89[4])
    defparam mode_160.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(n29194), .B(n29193), .C(mode), .D(n29303), .Z(n27480)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(76[18:71])
    defparam i1_4_lut.init = 16'h5554;
    
endmodule
//
// Verilog Description of module \shutter(DEV_ID=4,UART_ADDRESS_WIDTH=4) 
//

module \shutter(DEV_ID=4,UART_ADDRESS_WIDTH=4)  (\mode[1] , \mode[2] , n29224, 
            pin_io_out_44, \pin_intrpt[14] , pin_io_out_42, \pin_intrpt[12] , 
            reset_r, n1, \cs_decoded[8] , n2, pin_io_out_43, \pin_intrpt[13] , 
            mode, clk, clk_enable_169, n29239, \spi_data_r[0] ) /* synthesis syn_module_defined=1 */ ;
    input \mode[1] ;
    input \mode[2] ;
    output n29224;
    input pin_io_out_44;
    output \pin_intrpt[14] ;
    input pin_io_out_42;
    output \pin_intrpt[12] ;
    input reset_r;
    output n1;
    input \cs_decoded[8] ;
    output n2;
    input pin_io_out_43;
    output \pin_intrpt[13] ;
    output mode;
    input clk;
    input clk_enable_169;
    input n29239;
    input \spi_data_r[0] ;
    
    wire \pin_intrpt[14]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[14] */ ;   // c:/s_links/sources/mcm_top.v(102[46:56])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    LUT4 i22757_2_lut_rep_496 (.A(\mode[1] ), .B(\mode[2] ), .Z(n29224)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i22757_2_lut_rep_496.init = 16'h1111;
    LUT4 i4193_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(pin_io_out_44), 
         .Z(\pin_intrpt[14] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i4193_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_4106_i1_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(pin_io_out_42), 
         .Z(\pin_intrpt[12] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4106_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_3922_i1_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(reset_r), 
         .Z(n1)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_3922_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_3909_i2_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(\cs_decoded[8] ), 
         .Z(n2)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_3909_i2_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_4105_i1_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(pin_io_out_43), 
         .Z(\pin_intrpt[13] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4105_i1_2_lut_3_lut.init = 16'he0e0;
    FD1P3IX mode_160 (.D(\spi_data_r[0] ), .SP(clk_enable_169), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=508, LSE_RLINE=540 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(81[8] 89[4])
    defparam mode_160.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \io(DEV_ID=4,UART_ADDRESS_WIDTH=4) 
//

module \io(DEV_ID=4,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_166, 
            n29239, \spi_data_r[0] ) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_166;
    input n29239;
    input \spi_data_r[0] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    FD1P3IX mode_90 (.D(\spi_data_r[0] ), .SP(clk_enable_166), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=464, LSE_RLINE=496 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(80[8] 88[4])
    defparam mode_90.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \quad_decoder(DEV_ID=6) 
//

module \quad_decoder(DEV_ID=6)  (quad_count, clk_1MHz, \spi_data_out_r_39__N_2338[0] , 
            clk, \spi_data_out_r_39__N_2483[0] , \quad_b[6] , quad_buffer, 
            \pin_intrpt[20] , n29239, clk_enable_76, \spi_data_r[31] , 
            \spi_data_r[30] , \spi_data_r[29] , \spi_data_r[28] , \spi_data_r[27] , 
            \spi_data_r[26] , \spi_data_r[25] , \spi_data_r[24] , \spi_data_r[23] , 
            \spi_data_r[22] , \spi_data_r[21] , \spi_data_r[20] , \spi_data_r[19] , 
            \spi_data_r[0] , \spi_data_r[18] , \spi_data_r[17] , \spi_data_r[16] , 
            \spi_data_r[15] , \spi_data_r[14] , \spi_data_r[13] , \spi_data_r[12] , 
            \spi_data_r[11] , \spi_data_r[10] , \spi_data_r[9] , \spi_data_r[8] , 
            \spi_data_r[7] , \spi_data_r[6] , \spi_data_r[5] , \spi_data_r[4] , 
            \spi_data_r[3] , \spi_data_r[2] , \spi_data_r[1] , clk_enable_499, 
            n29762, resetn_c, GND_net, spi_data_out_r_39__N_2378, spi_data_out_r_39__N_2566, 
            quad_set_complete, \quad_a[6] , \spi_data_out_r_39__N_2338[31] , 
            \spi_data_out_r_39__N_2483[31] , \spi_data_out_r_39__N_2338[30] , 
            \spi_data_out_r_39__N_2483[30] , \spi_data_out_r_39__N_2338[29] , 
            \spi_data_out_r_39__N_2483[29] , \spi_data_out_r_39__N_2338[28] , 
            \spi_data_out_r_39__N_2483[28] , \spi_data_out_r_39__N_2338[27] , 
            \spi_data_out_r_39__N_2483[27] , \spi_data_out_r_39__N_2338[26] , 
            \spi_data_out_r_39__N_2483[26] , \spi_data_out_r_39__N_2338[25] , 
            \spi_data_out_r_39__N_2483[25] , \spi_data_out_r_39__N_2338[24] , 
            \spi_data_out_r_39__N_2483[24] , \spi_data_out_r_39__N_2338[23] , 
            \spi_data_out_r_39__N_2483[23] , \spi_data_out_r_39__N_2338[22] , 
            \spi_data_out_r_39__N_2483[22] , \spi_data_out_r_39__N_2338[21] , 
            \spi_data_out_r_39__N_2483[21] , \spi_data_out_r_39__N_2338[20] , 
            \spi_data_out_r_39__N_2483[20] , \spi_data_out_r_39__N_2338[19] , 
            \spi_data_out_r_39__N_2483[19] , \spi_data_out_r_39__N_2338[18] , 
            \spi_data_out_r_39__N_2483[18] , \spi_data_out_r_39__N_2338[17] , 
            \spi_data_out_r_39__N_2483[17] , \spi_data_out_r_39__N_2338[16] , 
            \spi_data_out_r_39__N_2483[16] , \spi_data_out_r_39__N_2338[15] , 
            \spi_data_out_r_39__N_2483[15] , \spi_data_out_r_39__N_2338[14] , 
            \spi_data_out_r_39__N_2483[14] , \spi_data_out_r_39__N_2338[13] , 
            \spi_data_out_r_39__N_2483[13] , \spi_data_out_r_39__N_2338[12] , 
            \spi_data_out_r_39__N_2483[12] , \spi_data_out_r_39__N_2338[11] , 
            \spi_data_out_r_39__N_2483[11] , \spi_data_out_r_39__N_2338[10] , 
            \spi_data_out_r_39__N_2483[10] , \spi_data_out_r_39__N_2338[9] , 
            \spi_data_out_r_39__N_2483[9] , \spi_data_out_r_39__N_2338[8] , 
            \spi_data_out_r_39__N_2483[8] , \spi_data_out_r_39__N_2338[7] , 
            \spi_data_out_r_39__N_2483[7] , \spi_data_out_r_39__N_2338[6] , 
            \spi_data_out_r_39__N_2483[6] , \spi_data_out_r_39__N_2338[5] , 
            \spi_data_out_r_39__N_2483[5] , \spi_data_out_r_39__N_2338[4] , 
            \spi_data_out_r_39__N_2483[4] , \spi_data_out_r_39__N_2338[3] , 
            \spi_data_out_r_39__N_2483[3] , \spi_data_out_r_39__N_2338[2] , 
            \spi_data_out_r_39__N_2483[2] , \spi_data_out_r_39__N_2338[1] , 
            \spi_data_out_r_39__N_2483[1] , pin_io_out_64, n29267, clk_enable_520, 
            n29092) /* synthesis syn_module_defined=1 */ ;
    output [31:0]quad_count;
    input clk_1MHz;
    output \spi_data_out_r_39__N_2338[0] ;
    input clk;
    input \spi_data_out_r_39__N_2483[0] ;
    input \quad_b[6] ;
    output [31:0]quad_buffer;
    input \pin_intrpt[20] ;
    input n29239;
    input clk_enable_76;
    input \spi_data_r[31] ;
    input \spi_data_r[30] ;
    input \spi_data_r[29] ;
    input \spi_data_r[28] ;
    input \spi_data_r[27] ;
    input \spi_data_r[26] ;
    input \spi_data_r[25] ;
    input \spi_data_r[24] ;
    input \spi_data_r[23] ;
    input \spi_data_r[22] ;
    input \spi_data_r[21] ;
    input \spi_data_r[20] ;
    input \spi_data_r[19] ;
    input \spi_data_r[0] ;
    input \spi_data_r[18] ;
    input \spi_data_r[17] ;
    input \spi_data_r[16] ;
    input \spi_data_r[15] ;
    input \spi_data_r[14] ;
    input \spi_data_r[13] ;
    input \spi_data_r[12] ;
    input \spi_data_r[11] ;
    input \spi_data_r[10] ;
    input \spi_data_r[9] ;
    input \spi_data_r[8] ;
    input \spi_data_r[7] ;
    input \spi_data_r[6] ;
    input \spi_data_r[5] ;
    input \spi_data_r[4] ;
    input \spi_data_r[3] ;
    input \spi_data_r[2] ;
    input \spi_data_r[1] ;
    input clk_enable_499;
    input n29762;
    input resetn_c;
    input GND_net;
    output spi_data_out_r_39__N_2378;
    input spi_data_out_r_39__N_2566;
    output quad_set_complete;
    input \quad_a[6] ;
    output \spi_data_out_r_39__N_2338[31] ;
    input \spi_data_out_r_39__N_2483[31] ;
    output \spi_data_out_r_39__N_2338[30] ;
    input \spi_data_out_r_39__N_2483[30] ;
    output \spi_data_out_r_39__N_2338[29] ;
    input \spi_data_out_r_39__N_2483[29] ;
    output \spi_data_out_r_39__N_2338[28] ;
    input \spi_data_out_r_39__N_2483[28] ;
    output \spi_data_out_r_39__N_2338[27] ;
    input \spi_data_out_r_39__N_2483[27] ;
    output \spi_data_out_r_39__N_2338[26] ;
    input \spi_data_out_r_39__N_2483[26] ;
    output \spi_data_out_r_39__N_2338[25] ;
    input \spi_data_out_r_39__N_2483[25] ;
    output \spi_data_out_r_39__N_2338[24] ;
    input \spi_data_out_r_39__N_2483[24] ;
    output \spi_data_out_r_39__N_2338[23] ;
    input \spi_data_out_r_39__N_2483[23] ;
    output \spi_data_out_r_39__N_2338[22] ;
    input \spi_data_out_r_39__N_2483[22] ;
    output \spi_data_out_r_39__N_2338[21] ;
    input \spi_data_out_r_39__N_2483[21] ;
    output \spi_data_out_r_39__N_2338[20] ;
    input \spi_data_out_r_39__N_2483[20] ;
    output \spi_data_out_r_39__N_2338[19] ;
    input \spi_data_out_r_39__N_2483[19] ;
    output \spi_data_out_r_39__N_2338[18] ;
    input \spi_data_out_r_39__N_2483[18] ;
    output \spi_data_out_r_39__N_2338[17] ;
    input \spi_data_out_r_39__N_2483[17] ;
    output \spi_data_out_r_39__N_2338[16] ;
    input \spi_data_out_r_39__N_2483[16] ;
    output \spi_data_out_r_39__N_2338[15] ;
    input \spi_data_out_r_39__N_2483[15] ;
    output \spi_data_out_r_39__N_2338[14] ;
    input \spi_data_out_r_39__N_2483[14] ;
    output \spi_data_out_r_39__N_2338[13] ;
    input \spi_data_out_r_39__N_2483[13] ;
    output \spi_data_out_r_39__N_2338[12] ;
    input \spi_data_out_r_39__N_2483[12] ;
    output \spi_data_out_r_39__N_2338[11] ;
    input \spi_data_out_r_39__N_2483[11] ;
    output \spi_data_out_r_39__N_2338[10] ;
    input \spi_data_out_r_39__N_2483[10] ;
    output \spi_data_out_r_39__N_2338[9] ;
    input \spi_data_out_r_39__N_2483[9] ;
    output \spi_data_out_r_39__N_2338[8] ;
    input \spi_data_out_r_39__N_2483[8] ;
    output \spi_data_out_r_39__N_2338[7] ;
    input \spi_data_out_r_39__N_2483[7] ;
    output \spi_data_out_r_39__N_2338[6] ;
    input \spi_data_out_r_39__N_2483[6] ;
    output \spi_data_out_r_39__N_2338[5] ;
    input \spi_data_out_r_39__N_2483[5] ;
    output \spi_data_out_r_39__N_2338[4] ;
    input \spi_data_out_r_39__N_2483[4] ;
    output \spi_data_out_r_39__N_2338[3] ;
    input \spi_data_out_r_39__N_2483[3] ;
    output \spi_data_out_r_39__N_2338[2] ;
    input \spi_data_out_r_39__N_2483[2] ;
    output \spi_data_out_r_39__N_2338[1] ;
    input \spi_data_out_r_39__N_2483[1] ;
    input pin_io_out_64;
    input n29267;
    input clk_enable_520;
    input n29092;
    
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire [1:0]sync /* synthesis ASYNC_REG="TRUE" */ ;   // c:/s_links/sources/quad_decoder.v(106[30:34])
    wire [1:0]AB /* synthesis ASYNC_REG="TRUE" */ ;   // c:/s_links/sources/quad_decoder.v(106[36:38])
    wire \pin_intrpt[20]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[20] */ ;   // c:/s_links/sources/mcm_top.v(102[46:56])
    
    wire clk_1MHz_enable_140, n26147;
    wire [3:0]n2471;
    
    wire n28552;
    wire [31:0]quad_set;   // c:/s_links/sources/quad_decoder.v(40[31:39])
    wire [1:0]quad_homing;   // c:/s_links/sources/quad_decoder.v(41[19:30])
    
    wire n25110, n11560;
    wire [31:0]n6431;
    
    wire n25109, n29003, n9480, n28952, n9471, n26745, n3, n27133, 
        n25823, n25825, n25841, n25839, n25861, n25859, n25881, 
        n6, n25879, n25901, quad_set_valid, n25899, n25921, n25919, 
        n25941, n25939, n25961, n25959, n25979, n25981, n26001, 
        n25999, n26021, n26019, n26041, n26039, n25108, n25107, 
        n25106, n25105, n25104, n25103, n25102, n25101, n25100, 
        n26073, n25099, n25098, n25097, n25096, n25095, n26071, 
        n26095, n26093, n26115, n26113, n26149, n26959, n13043, 
        n11446, n10, n4;
    
    FD1P3AX quad_count_i0_i0 (.D(n26147), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_2483[0] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX sync_i0 (.D(\quad_b[6] ), .CK(clk_1MHz), .Q(sync[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam sync_i0.GSR = "DISABLED";
    FD1S3AX AB_i0 (.D(sync[0]), .CK(clk_1MHz), .Q(AB[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam AB_i0.GSR = "DISABLED";
    FD1S3AX quad_buffer_i0 (.D(quad_count[0]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i0.GSR = "DISABLED";
    FD1S3JX state_FSM_i0 (.D(n28552), .CK(clk_1MHz), .PD(n29239), .Q(n2471[0]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i0.GSR = "DISABLED";
    FD1P3IX quad_set__i31 (.D(\spi_data_r[31] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i31.GSR = "DISABLED";
    FD1P3IX quad_set__i30 (.D(\spi_data_r[30] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i30.GSR = "DISABLED";
    FD1P3IX quad_set__i29 (.D(\spi_data_r[29] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i29.GSR = "DISABLED";
    FD1P3IX quad_set__i28 (.D(\spi_data_r[28] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i28.GSR = "DISABLED";
    FD1P3IX quad_set__i27 (.D(\spi_data_r[27] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i27.GSR = "DISABLED";
    FD1P3IX quad_set__i26 (.D(\spi_data_r[26] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i26.GSR = "DISABLED";
    FD1P3IX quad_set__i25 (.D(\spi_data_r[25] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i25.GSR = "DISABLED";
    FD1P3IX quad_set__i24 (.D(\spi_data_r[24] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i24.GSR = "DISABLED";
    FD1P3IX quad_set__i23 (.D(\spi_data_r[23] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i23.GSR = "DISABLED";
    FD1P3IX quad_set__i22 (.D(\spi_data_r[22] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i22.GSR = "DISABLED";
    FD1P3IX quad_set__i21 (.D(\spi_data_r[21] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i21.GSR = "DISABLED";
    FD1P3IX quad_set__i20 (.D(\spi_data_r[20] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i20.GSR = "DISABLED";
    FD1P3IX quad_set__i19 (.D(\spi_data_r[19] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i19.GSR = "DISABLED";
    FD1P3IX quad_set__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i0.GSR = "DISABLED";
    FD1P3IX quad_set__i18 (.D(\spi_data_r[18] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i18.GSR = "DISABLED";
    FD1P3IX quad_set__i17 (.D(\spi_data_r[17] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i17.GSR = "DISABLED";
    FD1P3IX quad_set__i16 (.D(\spi_data_r[16] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i16.GSR = "DISABLED";
    FD1P3IX quad_set__i15 (.D(\spi_data_r[15] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i15.GSR = "DISABLED";
    FD1P3IX quad_set__i14 (.D(\spi_data_r[14] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i14.GSR = "DISABLED";
    FD1P3IX quad_set__i13 (.D(\spi_data_r[13] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i13.GSR = "DISABLED";
    FD1P3IX quad_set__i12 (.D(\spi_data_r[12] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i12.GSR = "DISABLED";
    FD1P3IX quad_set__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i11.GSR = "DISABLED";
    FD1P3IX quad_set__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i10.GSR = "DISABLED";
    FD1P3IX quad_set__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i9.GSR = "DISABLED";
    FD1P3IX quad_set__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i8.GSR = "DISABLED";
    FD1P3IX quad_set__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i7.GSR = "DISABLED";
    FD1P3IX quad_set__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i6.GSR = "DISABLED";
    FD1P3IX quad_set__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i5.GSR = "DISABLED";
    FD1P3IX quad_set__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i4.GSR = "DISABLED";
    FD1P3IX quad_set__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i3.GSR = "DISABLED";
    FD1P3IX quad_set__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i2.GSR = "DISABLED";
    FD1P3IX quad_set__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_76), .CD(n29239), 
            .CK(clk), .Q(quad_set[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i1.GSR = "DISABLED";
    FD1P3IX quad_homing__i0 (.D(n29762), .SP(clk_enable_499), .CD(n29239), 
            .CK(clk), .Q(quad_homing[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam quad_homing__i0.GSR = "DISABLED";
    CCU2D add_2112_33 (.A0(resetn_c), .B0(n11560), .C0(quad_count[30]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[31]), 
          .D1(GND_net), .CIN(n25110), .S0(n6431[30]), .S1(n6431[31]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_33.INIT0 = 16'hd2d2;
    defparam add_2112_33.INIT1 = 16'hd2d2;
    defparam add_2112_33.INJECT1_0 = "NO";
    defparam add_2112_33.INJECT1_1 = "NO";
    CCU2D add_2112_31 (.A0(resetn_c), .B0(n11560), .C0(quad_count[28]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[29]), 
          .D1(GND_net), .CIN(n25109), .COUT(n25110), .S0(n6431[28]), 
          .S1(n6431[29]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_31.INIT0 = 16'hd2d2;
    defparam add_2112_31.INIT1 = 16'hd2d2;
    defparam add_2112_31.INJECT1_0 = "NO";
    defparam add_2112_31.INJECT1_1 = "NO";
    FD1S3IX state_FSM_i3 (.D(n29003), .CK(clk_1MHz), .CD(n29239), .Q(n2471[3]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i3.GSR = "DISABLED";
    FD1S3IX state_FSM_i2 (.D(n9480), .CK(clk_1MHz), .CD(n29239), .Q(n2471[2]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i2.GSR = "DISABLED";
    FD1S3IX state_FSM_i1 (.D(n28952), .CK(clk_1MHz), .CD(n29239), .Q(n2471[1]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i1.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut (.A(n2471[3]), .B(AB[0]), .C(AB[1]), .D(n9471), 
         .Z(n26745)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i1_4_lut_4_lut.init = 16'h96c3;
    LUT4 i31_4_lut (.A(n6431[31]), .B(quad_set[31]), .C(n3), .D(n27133), 
         .Z(n25823)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut.init = 16'hcac0;
    LUT4 i31_4_lut_adj_971 (.A(n6431[30]), .B(quad_set[30]), .C(n3), .D(n27133), 
         .Z(n25825)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_971.init = 16'hcac0;
    LUT4 i31_4_lut_adj_972 (.A(n6431[29]), .B(quad_set[29]), .C(n3), .D(n27133), 
         .Z(n25841)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_972.init = 16'hcac0;
    LUT4 i31_4_lut_adj_973 (.A(n6431[28]), .B(quad_set[28]), .C(n3), .D(n27133), 
         .Z(n25839)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_973.init = 16'hcac0;
    LUT4 i31_4_lut_adj_974 (.A(n6431[27]), .B(quad_set[27]), .C(n3), .D(n27133), 
         .Z(n25861)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_974.init = 16'hcac0;
    LUT4 i31_4_lut_adj_975 (.A(n6431[26]), .B(quad_set[26]), .C(n3), .D(n27133), 
         .Z(n25859)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_975.init = 16'hcac0;
    LUT4 i31_4_lut_adj_976 (.A(n6431[25]), .B(quad_set[25]), .C(n3), .D(n27133), 
         .Z(n25881)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_976.init = 16'hcac0;
    LUT4 i4706_4_lut_4_lut (.A(n2471[2]), .B(AB[0]), .C(AB[1]), .D(n6), 
         .Z(n9480)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C (D))))) */ ;   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam i4706_4_lut_4_lut.init = 16'h3828;
    LUT4 i31_4_lut_adj_977 (.A(n6431[24]), .B(quad_set[24]), .C(n3), .D(n27133), 
         .Z(n25879)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_977.init = 16'hcac0;
    LUT4 i31_4_lut_adj_978 (.A(n6431[23]), .B(quad_set[23]), .C(n3), .D(n27133), 
         .Z(n25901)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_978.init = 16'hcac0;
    FD1S3IX i41_407 (.D(spi_data_out_r_39__N_2566), .CK(clk), .CD(n29239), 
            .Q(spi_data_out_r_39__N_2378)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam i41_407.GSR = "DISABLED";
    FD1S3IX quad_set_complete_451 (.D(quad_set_valid), .CK(clk_1MHz), .CD(n29239), 
            .Q(quad_set_complete)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_set_complete_451.GSR = "DISABLED";
    LUT4 i31_4_lut_adj_979 (.A(n6431[22]), .B(quad_set[22]), .C(n3), .D(n27133), 
         .Z(n25899)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_979.init = 16'hcac0;
    LUT4 i31_4_lut_adj_980 (.A(n6431[21]), .B(quad_set[21]), .C(n3), .D(n27133), 
         .Z(n25921)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_980.init = 16'hcac0;
    LUT4 i31_4_lut_adj_981 (.A(n6431[20]), .B(quad_set[20]), .C(n3), .D(n27133), 
         .Z(n25919)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_981.init = 16'hcac0;
    LUT4 i31_4_lut_adj_982 (.A(n6431[19]), .B(quad_set[19]), .C(n3), .D(n27133), 
         .Z(n25941)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_982.init = 16'hcac0;
    LUT4 i31_4_lut_adj_983 (.A(n6431[18]), .B(quad_set[18]), .C(n3), .D(n27133), 
         .Z(n25939)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_983.init = 16'hcac0;
    LUT4 i31_4_lut_adj_984 (.A(n6431[17]), .B(quad_set[17]), .C(n3), .D(n27133), 
         .Z(n25961)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_984.init = 16'hcac0;
    LUT4 i31_4_lut_adj_985 (.A(n6431[16]), .B(quad_set[16]), .C(n3), .D(n27133), 
         .Z(n25959)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_985.init = 16'hcac0;
    LUT4 n6_bdd_4_lut (.A(n6), .B(n2471[1]), .C(AB[0]), .D(AB[1]), .Z(n28952)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C (D)+!C !(D))+!B))) */ ;
    defparam n6_bdd_4_lut.init = 16'h0ce0;
    LUT4 i1_2_lut (.A(n2471[0]), .B(n2471[3]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i31_4_lut_adj_986 (.A(n6431[15]), .B(quad_set[15]), .C(n3), .D(n27133), 
         .Z(n25979)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_986.init = 16'hcac0;
    LUT4 i31_4_lut_adj_987 (.A(n6431[14]), .B(quad_set[14]), .C(n3), .D(n27133), 
         .Z(n25981)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_987.init = 16'hcac0;
    LUT4 i31_4_lut_adj_988 (.A(n6431[13]), .B(quad_set[13]), .C(n3), .D(n27133), 
         .Z(n26001)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_988.init = 16'hcac0;
    LUT4 AB_1__bdd_4_lut (.A(AB[1]), .B(n2471[3]), .C(AB[0]), .D(n9471), 
         .Z(n29003)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam AB_1__bdd_4_lut.init = 16'ha484;
    LUT4 i31_4_lut_adj_989 (.A(n6431[12]), .B(quad_set[12]), .C(n3), .D(n27133), 
         .Z(n25999)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_989.init = 16'hcac0;
    LUT4 i31_4_lut_adj_990 (.A(n6431[11]), .B(quad_set[11]), .C(n3), .D(n27133), 
         .Z(n26021)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_990.init = 16'hcac0;
    LUT4 AB_1__bdd_4_lut_23135 (.A(AB[1]), .B(n2471[0]), .C(AB[0]), .D(n9471), 
         .Z(n28552)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B (C+!(D)))) */ ;
    defparam AB_1__bdd_4_lut_23135.init = 16'h8584;
    LUT4 i31_4_lut_adj_991 (.A(n6431[10]), .B(quad_set[10]), .C(n3), .D(n27133), 
         .Z(n26019)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_991.init = 16'hcac0;
    LUT4 i31_4_lut_adj_992 (.A(n6431[9]), .B(quad_set[9]), .C(n3), .D(n27133), 
         .Z(n26041)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_992.init = 16'hcac0;
    LUT4 i31_4_lut_adj_993 (.A(n6431[8]), .B(quad_set[8]), .C(n3), .D(n27133), 
         .Z(n26039)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_993.init = 16'hcac0;
    FD1S3AX quad_buffer_i31 (.D(quad_count[31]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i31.GSR = "DISABLED";
    FD1S3AX quad_buffer_i30 (.D(quad_count[30]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i30.GSR = "DISABLED";
    FD1S3AX quad_buffer_i29 (.D(quad_count[29]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i29.GSR = "DISABLED";
    FD1S3AX quad_buffer_i28 (.D(quad_count[28]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i28.GSR = "DISABLED";
    FD1S3AX quad_buffer_i27 (.D(quad_count[27]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i27.GSR = "DISABLED";
    FD1S3AX quad_buffer_i26 (.D(quad_count[26]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i26.GSR = "DISABLED";
    FD1S3AX quad_buffer_i25 (.D(quad_count[25]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i25.GSR = "DISABLED";
    FD1S3AX quad_buffer_i24 (.D(quad_count[24]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i24.GSR = "DISABLED";
    FD1S3AX quad_buffer_i23 (.D(quad_count[23]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i23.GSR = "DISABLED";
    CCU2D add_2112_29 (.A0(resetn_c), .B0(n11560), .C0(quad_count[26]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[27]), 
          .D1(GND_net), .CIN(n25108), .COUT(n25109), .S0(n6431[26]), 
          .S1(n6431[27]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_29.INIT0 = 16'hd2d2;
    defparam add_2112_29.INIT1 = 16'hd2d2;
    defparam add_2112_29.INJECT1_0 = "NO";
    defparam add_2112_29.INJECT1_1 = "NO";
    FD1S3AX quad_buffer_i22 (.D(quad_count[22]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i22.GSR = "DISABLED";
    FD1S3AX quad_buffer_i21 (.D(quad_count[21]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i21.GSR = "DISABLED";
    FD1S3AX quad_buffer_i20 (.D(quad_count[20]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i20.GSR = "DISABLED";
    FD1S3AX quad_buffer_i19 (.D(quad_count[19]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i19.GSR = "DISABLED";
    FD1S3AX quad_buffer_i18 (.D(quad_count[18]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i18.GSR = "DISABLED";
    FD1S3AX quad_buffer_i17 (.D(quad_count[17]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i17.GSR = "DISABLED";
    FD1S3AX quad_buffer_i16 (.D(quad_count[16]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i16.GSR = "DISABLED";
    FD1S3AX quad_buffer_i15 (.D(quad_count[15]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i15.GSR = "DISABLED";
    FD1S3AX quad_buffer_i14 (.D(quad_count[14]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i14.GSR = "DISABLED";
    FD1S3AX quad_buffer_i13 (.D(quad_count[13]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i13.GSR = "DISABLED";
    FD1S3AX quad_buffer_i12 (.D(quad_count[12]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i12.GSR = "DISABLED";
    FD1S3AX quad_buffer_i11 (.D(quad_count[11]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i11.GSR = "DISABLED";
    FD1S3AX quad_buffer_i10 (.D(quad_count[10]), .CK(\pin_intrpt[20] ), 
            .Q(quad_buffer[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i10.GSR = "DISABLED";
    FD1S3AX quad_buffer_i9 (.D(quad_count[9]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i9.GSR = "DISABLED";
    FD1S3AX quad_buffer_i8 (.D(quad_count[8]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i8.GSR = "DISABLED";
    FD1S3AX quad_buffer_i7 (.D(quad_count[7]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i7.GSR = "DISABLED";
    FD1S3AX quad_buffer_i6 (.D(quad_count[6]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i6.GSR = "DISABLED";
    FD1S3AX quad_buffer_i5 (.D(quad_count[5]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i5.GSR = "DISABLED";
    FD1S3AX quad_buffer_i4 (.D(quad_count[4]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i4.GSR = "DISABLED";
    FD1S3AX quad_buffer_i3 (.D(quad_count[3]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i3.GSR = "DISABLED";
    FD1S3AX quad_buffer_i2 (.D(quad_count[2]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i2.GSR = "DISABLED";
    FD1S3AX quad_buffer_i1 (.D(quad_count[1]), .CK(\pin_intrpt[20] ), .Q(quad_buffer[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i1.GSR = "DISABLED";
    FD1S3AX AB_i1 (.D(sync[1]), .CK(clk_1MHz), .Q(AB[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam AB_i1.GSR = "DISABLED";
    FD1S3AX sync_i1 (.D(\quad_a[6] ), .CK(clk_1MHz), .Q(sync[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam sync_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_2483[31] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i31 (.D(\spi_data_out_r_39__N_2483[30] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i30 (.D(\spi_data_out_r_39__N_2483[29] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i29 (.D(\spi_data_out_r_39__N_2483[28] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i28 (.D(\spi_data_out_r_39__N_2483[27] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i27 (.D(\spi_data_out_r_39__N_2483[26] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i26 (.D(\spi_data_out_r_39__N_2483[25] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i25 (.D(\spi_data_out_r_39__N_2483[24] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i24 (.D(\spi_data_out_r_39__N_2483[23] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i23 (.D(\spi_data_out_r_39__N_2483[22] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i22 (.D(\spi_data_out_r_39__N_2483[21] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i21 (.D(\spi_data_out_r_39__N_2483[20] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i20 (.D(\spi_data_out_r_39__N_2483[19] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i19 (.D(\spi_data_out_r_39__N_2483[18] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i18 (.D(\spi_data_out_r_39__N_2483[17] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i17 (.D(\spi_data_out_r_39__N_2483[16] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i16 (.D(\spi_data_out_r_39__N_2483[15] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_2483[14] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_2483[13] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_2483[12] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_2483[11] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_2483[10] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_2483[9] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_2483[8] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_2483[7] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_2483[6] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_2483[5] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_2483[4] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_2483[3] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_2483[2] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_2483[1] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2338[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    CCU2D add_2112_27 (.A0(resetn_c), .B0(n11560), .C0(quad_count[24]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[25]), 
          .D1(GND_net), .CIN(n25107), .COUT(n25108), .S0(n6431[24]), 
          .S1(n6431[25]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_27.INIT0 = 16'hd2d2;
    defparam add_2112_27.INIT1 = 16'hd2d2;
    defparam add_2112_27.INJECT1_0 = "NO";
    defparam add_2112_27.INJECT1_1 = "NO";
    CCU2D add_2112_25 (.A0(resetn_c), .B0(n11560), .C0(quad_count[22]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[23]), 
          .D1(GND_net), .CIN(n25106), .COUT(n25107), .S0(n6431[22]), 
          .S1(n6431[23]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_25.INIT0 = 16'hd2d2;
    defparam add_2112_25.INIT1 = 16'hd2d2;
    defparam add_2112_25.INJECT1_0 = "NO";
    defparam add_2112_25.INJECT1_1 = "NO";
    CCU2D add_2112_23 (.A0(resetn_c), .B0(n11560), .C0(quad_count[20]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[21]), 
          .D1(GND_net), .CIN(n25105), .COUT(n25106), .S0(n6431[20]), 
          .S1(n6431[21]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_23.INIT0 = 16'hd2d2;
    defparam add_2112_23.INIT1 = 16'hd2d2;
    defparam add_2112_23.INJECT1_0 = "NO";
    defparam add_2112_23.INJECT1_1 = "NO";
    CCU2D add_2112_21 (.A0(resetn_c), .B0(n11560), .C0(quad_count[18]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[19]), 
          .D1(GND_net), .CIN(n25104), .COUT(n25105), .S0(n6431[18]), 
          .S1(n6431[19]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_21.INIT0 = 16'hd2d2;
    defparam add_2112_21.INIT1 = 16'hd2d2;
    defparam add_2112_21.INJECT1_0 = "NO";
    defparam add_2112_21.INJECT1_1 = "NO";
    CCU2D add_2112_19 (.A0(resetn_c), .B0(n11560), .C0(quad_count[16]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[17]), 
          .D1(GND_net), .CIN(n25103), .COUT(n25104), .S0(n6431[16]), 
          .S1(n6431[17]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_19.INIT0 = 16'hd2d2;
    defparam add_2112_19.INIT1 = 16'hd2d2;
    defparam add_2112_19.INJECT1_0 = "NO";
    defparam add_2112_19.INJECT1_1 = "NO";
    CCU2D add_2112_17 (.A0(resetn_c), .B0(n11560), .C0(quad_count[14]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[15]), 
          .D1(GND_net), .CIN(n25102), .COUT(n25103), .S0(n6431[14]), 
          .S1(n6431[15]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_17.INIT0 = 16'hd2d2;
    defparam add_2112_17.INIT1 = 16'hd2d2;
    defparam add_2112_17.INJECT1_0 = "NO";
    defparam add_2112_17.INJECT1_1 = "NO";
    CCU2D add_2112_15 (.A0(resetn_c), .B0(n11560), .C0(quad_count[12]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[13]), 
          .D1(GND_net), .CIN(n25101), .COUT(n25102), .S0(n6431[12]), 
          .S1(n6431[13]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_15.INIT0 = 16'hd2d2;
    defparam add_2112_15.INIT1 = 16'hd2d2;
    defparam add_2112_15.INJECT1_0 = "NO";
    defparam add_2112_15.INJECT1_1 = "NO";
    CCU2D add_2112_13 (.A0(resetn_c), .B0(n11560), .C0(quad_count[10]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[11]), 
          .D1(GND_net), .CIN(n25100), .COUT(n25101), .S0(n6431[10]), 
          .S1(n6431[11]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_13.INIT0 = 16'hd2d2;
    defparam add_2112_13.INIT1 = 16'hd2d2;
    defparam add_2112_13.INJECT1_0 = "NO";
    defparam add_2112_13.INJECT1_1 = "NO";
    LUT4 i31_4_lut_adj_994 (.A(n6431[7]), .B(quad_set[7]), .C(n3), .D(n27133), 
         .Z(n26073)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_994.init = 16'hcac0;
    CCU2D add_2112_11 (.A0(resetn_c), .B0(n11560), .C0(quad_count[8]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[9]), 
          .D1(GND_net), .CIN(n25099), .COUT(n25100), .S0(n6431[8]), 
          .S1(n6431[9]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_11.INIT0 = 16'hd2d2;
    defparam add_2112_11.INIT1 = 16'hd2d2;
    defparam add_2112_11.INJECT1_0 = "NO";
    defparam add_2112_11.INJECT1_1 = "NO";
    CCU2D add_2112_9 (.A0(resetn_c), .B0(n11560), .C0(quad_count[6]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[7]), 
          .D1(GND_net), .CIN(n25098), .COUT(n25099), .S0(n6431[6]), 
          .S1(n6431[7]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_9.INIT0 = 16'hd2d2;
    defparam add_2112_9.INIT1 = 16'hd2d2;
    defparam add_2112_9.INJECT1_0 = "NO";
    defparam add_2112_9.INJECT1_1 = "NO";
    CCU2D add_2112_7 (.A0(resetn_c), .B0(n11560), .C0(quad_count[4]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[5]), 
          .D1(GND_net), .CIN(n25097), .COUT(n25098), .S0(n6431[4]), 
          .S1(n6431[5]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_7.INIT0 = 16'hd2d2;
    defparam add_2112_7.INIT1 = 16'hd2d2;
    defparam add_2112_7.INJECT1_0 = "NO";
    defparam add_2112_7.INJECT1_1 = "NO";
    CCU2D add_2112_5 (.A0(resetn_c), .B0(n11560), .C0(quad_count[2]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[3]), 
          .D1(GND_net), .CIN(n25096), .COUT(n25097), .S0(n6431[2]), 
          .S1(n6431[3]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_5.INIT0 = 16'hd2d2;
    defparam add_2112_5.INIT1 = 16'hd2d2;
    defparam add_2112_5.INJECT1_0 = "NO";
    defparam add_2112_5.INJECT1_1 = "NO";
    CCU2D add_2112_3 (.A0(resetn_c), .B0(n11560), .C0(quad_count[0]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11560), .C1(quad_count[1]), 
          .D1(GND_net), .CIN(n25095), .COUT(n25096), .S0(n6431[0]), 
          .S1(n6431[1]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_3.INIT0 = 16'h2d2d;
    defparam add_2112_3.INIT1 = 16'hd2d2;
    defparam add_2112_3.INJECT1_0 = "NO";
    defparam add_2112_3.INJECT1_1 = "NO";
    CCU2D add_2112_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(resetn_c), .B1(n11560), .C1(GND_net), .D1(GND_net), .COUT(n25095));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2112_1.INIT0 = 16'hF000;
    defparam add_2112_1.INIT1 = 16'hdddd;
    defparam add_2112_1.INJECT1_0 = "NO";
    defparam add_2112_1.INJECT1_1 = "NO";
    LUT4 i31_4_lut_adj_995 (.A(n6431[6]), .B(quad_set[6]), .C(n3), .D(n27133), 
         .Z(n26071)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_995.init = 16'hcac0;
    LUT4 i31_4_lut_adj_996 (.A(n6431[5]), .B(quad_set[5]), .C(n3), .D(n27133), 
         .Z(n26095)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_996.init = 16'hcac0;
    LUT4 i31_4_lut_adj_997 (.A(n6431[4]), .B(quad_set[4]), .C(n3), .D(n27133), 
         .Z(n26093)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_997.init = 16'hcac0;
    LUT4 i31_4_lut_adj_998 (.A(n6431[3]), .B(quad_set[3]), .C(n3), .D(n27133), 
         .Z(n26115)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_998.init = 16'hcac0;
    LUT4 i31_4_lut_adj_999 (.A(n6431[2]), .B(quad_set[2]), .C(n3), .D(n27133), 
         .Z(n26113)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_999.init = 16'hcac0;
    LUT4 i31_4_lut_adj_1000 (.A(n6431[1]), .B(quad_set[1]), .C(n3), .D(n27133), 
         .Z(n26149)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_1000.init = 16'hcac0;
    FD1P3AX quad_count_i0_i31 (.D(n25823), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i31.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i30 (.D(n25825), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i30.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i29 (.D(n25841), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i29.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i28 (.D(n25839), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i28.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i27 (.D(n25861), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i27.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i26 (.D(n25859), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i26.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i25 (.D(n25881), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i25.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i24 (.D(n25879), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i24.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i23 (.D(n25901), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i23.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i22 (.D(n25899), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i22.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i21 (.D(n25921), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i21.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i20 (.D(n25919), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i20.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i19 (.D(n25941), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i19.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i18 (.D(n25939), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i18.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i17 (.D(n25961), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i17.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i16 (.D(n25959), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i16.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i15 (.D(n25979), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i15.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i14 (.D(n25981), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i14.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i13 (.D(n26001), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i13.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i12 (.D(n25999), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i12.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i11 (.D(n26021), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i11.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i10 (.D(n26019), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i10.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i9 (.D(n26041), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i9.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i8 (.D(n26039), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i8.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i7 (.D(n26073), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i7.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i6 (.D(n26071), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i6.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i5 (.D(n26095), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i5.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i4 (.D(n26093), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i4.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i3 (.D(n26115), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i3.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i2 (.D(n26113), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i1 (.D(n26149), .SP(clk_1MHz_enable_140), .CK(clk_1MHz), 
            .Q(quad_count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i1.GSR = "DISABLED";
    LUT4 i2_3_lut_4_lut (.A(quad_homing[0]), .B(pin_io_out_64), .C(n29267), 
         .D(quad_homing[1]), .Z(n26959)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfff7;
    LUT4 i3_3_lut_4_lut (.A(quad_homing[0]), .B(pin_io_out_64), .C(n29267), 
         .D(quad_homing[1]), .Z(n13043)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i3_3_lut_4_lut.init = 16'h0008;
    LUT4 i5150_3_lut_4_lut (.A(AB[0]), .B(AB[1]), .C(n2471[3]), .D(n11446), 
         .Z(n11560)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // c:/s_links/sources/quad_decoder.v(162[19:30])
    defparam i5150_3_lut_4_lut.init = 16'hbfb0;
    FD1P3IX quad_homing__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_499), .CD(n29239), 
            .CK(clk), .Q(quad_homing[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam quad_homing__i1.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(n2471[1]), .B(n10), .C(n2471[2]), .D(n2471[3]), 
         .Z(n4)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i1_4_lut.init = 16'h33c9;
    LUT4 reduce_or_662_i1_2_lut (.A(n2471[2]), .B(n2471[1]), .Z(n9471)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam reduce_or_662_i1_2_lut.init = 16'heeee;
    LUT4 i15_2_lut (.A(AB[1]), .B(AB[0]), .Z(n10)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(155[16] 158[10])
    defparam i15_2_lut.init = 16'h6666;
    FD1P3IX quad_set_valid_404 (.D(n29092), .SP(clk_enable_520), .CD(n29239), 
            .CK(clk), .Q(quad_set_valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set_valid_404.GSR = "DISABLED";
    LUT4 i5149_4_lut (.A(AB[0]), .B(AB[1]), .C(n2471[2]), .D(n2471[1]), 
         .Z(n11446)) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A (B+!(C))) */ ;
    defparam i5149_4_lut.init = 16'he7ed;
    LUT4 i22855_4_lut (.A(n26745), .B(resetn_c), .C(quad_set_valid), .D(n13043), 
         .Z(clk_1MHz_enable_140)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i22855_4_lut.init = 16'hfff7;
    LUT4 i31_4_lut_adj_1001 (.A(n6431[0]), .B(quad_set[0]), .C(n3), .D(n27133), 
         .Z(n26147)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_1001.init = 16'hcac0;
    LUT4 i2_4_lut (.A(n26959), .B(quad_set_valid), .C(n4), .D(resetn_c), 
         .Z(n3)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'h8000;
    LUT4 i1_3_lut (.A(resetn_c), .B(n13043), .C(n4), .Z(n27133)) /* synthesis lut_function=(!((B (C))+!A)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i1_3_lut.init = 16'h2a2a;
    
endmodule
//
// Verilog Description of module \io(DEV_ID=5,UART_ADDRESS_WIDTH=4) 
//

module \io(DEV_ID=5,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_182, 
            n29239, \spi_data_r[0] ) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_182;
    input n29239;
    input \spi_data_r[0] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    FD1P3IX mode_90 (.D(\spi_data_r[0] ), .SP(clk_enable_182), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=464, LSE_RLINE=496 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(80[8] 88[4])
    defparam mode_90.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \io(UART_ADDRESS_WIDTH=4) 
//

module \io(UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_167, n29239, 
            \spi_data_r[0] , \spi_cmd_r[2] , \spi_addr_r[2] , n29256, 
            n29101, resetn_c, clk_enable_178, n19233, \spi_addr_r[0] , 
            \spi_cmd_r[1] , n29288, n65, n29110, \spi_cmd_r[0] , n27058, 
            n13074, n29213, \spi_cmd[1] , \spi_addr_r[3] , spi_sdo_valid_N_297, 
            spi_sdo_valid_N_296, \spi_cmd[2] , \spi_cmd[15] , n29761, 
            n19084, n27618, n31, \spi_cmd[4] , n29144, n29182, n29169, 
            n29114, \spi_addr_r[1] , n29214, n29105, n29211, n27225, 
            n29120) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_167;
    input n29239;
    input \spi_data_r[0] ;
    input \spi_cmd_r[2] ;
    input \spi_addr_r[2] ;
    output n29256;
    input n29101;
    input resetn_c;
    output clk_enable_178;
    output n19233;
    input \spi_addr_r[0] ;
    input \spi_cmd_r[1] ;
    output n29288;
    input n65;
    output n29110;
    input \spi_cmd_r[0] ;
    output n27058;
    output n13074;
    output n29213;
    input \spi_cmd[1] ;
    input \spi_addr_r[3] ;
    output spi_sdo_valid_N_297;
    input spi_sdo_valid_N_296;
    input \spi_cmd[2] ;
    input \spi_cmd[15] ;
    input n29761;
    input n19084;
    input n27618;
    input n31;
    input \spi_cmd[4] ;
    input n29144;
    input n29182;
    input n29169;
    output n29114;
    input \spi_addr_r[1] ;
    input n29214;
    output n29105;
    input n29211;
    input n27225;
    output n29120;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    wire n13, n27653;
    
    FD1P3IX mode_90 (.D(\spi_data_r[0] ), .SP(clk_enable_167), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=464, LSE_RLINE=496 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(80[8] 88[4])
    defparam mode_90.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_528 (.A(\spi_cmd_r[2] ), .B(\spi_addr_r[2] ), .Z(n29256)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/s_links/sources/slot_cards/slider_io.v(83[15:49])
    defparam i1_2_lut_rep_528.init = 16'h4444;
    LUT4 i1_3_lut_3_lut_4_lut (.A(\spi_cmd_r[2] ), .B(\spi_addr_r[2] ), 
         .C(n29101), .D(resetn_c), .Z(clk_enable_178)) /* synthesis lut_function=(!(A (D)+!A !(B (C+!(D))+!B !(D)))) */ ;   // c:/s_links/sources/slot_cards/slider_io.v(83[15:49])
    defparam i1_3_lut_3_lut_4_lut.init = 16'h40ff;
    LUT4 i14306_2_lut (.A(\spi_cmd_r[2] ), .B(\spi_addr_r[2] ), .Z(n19233)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14306_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_rep_560 (.A(\spi_addr_r[0] ), .B(\spi_cmd_r[1] ), .Z(n29288)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_560.init = 16'h2222;
    LUT4 i2_3_lut_rep_382_4_lut (.A(\spi_addr_r[0] ), .B(\spi_cmd_r[1] ), 
         .C(n65), .D(n19233), .Z(n29110)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i2_3_lut_rep_382_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\spi_cmd_r[0] ), .B(\spi_cmd_r[1] ), .C(\spi_cmd_r[2] ), 
         .D(\spi_addr_r[0] ), .Z(n27058)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_3_lut (.A(\spi_cmd_r[0] ), .B(\spi_cmd_r[1] ), .C(\spi_addr_r[0] ), 
         .Z(n13074)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h0202;
    LUT4 i1_2_lut_rep_485_3_lut (.A(\spi_cmd_r[0] ), .B(\spi_cmd_r[1] ), 
         .C(\spi_addr_r[0] ), .Z(n29213)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_rep_485_3_lut.init = 16'h2020;
    LUT4 i7_4_lut (.A(n13), .B(\spi_cmd[1] ), .C(n27653), .D(\spi_addr_r[3] ), 
         .Z(spi_sdo_valid_N_297)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i7_4_lut.init = 16'h0200;
    LUT4 i5_4_lut (.A(spi_sdo_valid_N_296), .B(\spi_cmd[2] ), .C(\spi_cmd[15] ), 
         .D(n29761), .Z(n13)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i5_4_lut.init = 16'h2000;
    LUT4 i22481_4_lut (.A(n19084), .B(n27618), .C(n31), .D(\spi_cmd[4] ), 
         .Z(n27653)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22481_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_386_3_lut_4_lut (.A(\spi_cmd_r[2] ), .B(n29144), .C(n29182), 
         .D(n29169), .Z(n29114)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/s_links/sources/slot_cards/slider_io.v(83[15:49])
    defparam i1_2_lut_rep_386_3_lut_4_lut.init = 16'h0004;
    LUT4 i1_2_lut_rep_377_3_lut_4_lut (.A(\spi_cmd_r[2] ), .B(n29144), .C(\spi_addr_r[1] ), 
         .D(n29214), .Z(n29105)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/s_links/sources/slot_cards/slider_io.v(83[15:49])
    defparam i1_2_lut_rep_377_3_lut_4_lut.init = 16'h0004;
    LUT4 i2_3_lut_rep_392_4_lut (.A(\spi_cmd_r[2] ), .B(n29144), .C(n29211), 
         .D(n27225), .Z(n29120)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/s_links/sources/slot_cards/slider_io.v(83[15:49])
    defparam i2_3_lut_rep_392_4_lut.init = 16'h4000;
    
endmodule
//
// Verilog Description of module \io(DEV_ID=2,UART_ADDRESS_WIDTH=4) 
//

module \io(DEV_ID=2,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_202, 
            n29239, \spi_data_r[0] ) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_202;
    input n29239;
    input \spi_data_r[0] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    FD1P3IX mode_90 (.D(\spi_data_r[0] ), .SP(clk_enable_202), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=464, LSE_RLINE=496 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(80[8] 88[4])
    defparam mode_90.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \io(DEV_ID=1,UART_ADDRESS_WIDTH=4) 
//

module \io(DEV_ID=1,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_197, 
            n29239, \spi_data_r[0] ) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_197;
    input n29239;
    input \spi_data_r[0] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    FD1P3IX mode_90 (.D(\spi_data_r[0] ), .SP(clk_enable_197), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=464, LSE_RLINE=496 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(80[8] 88[4])
    defparam mode_90.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \servo(DEV_ID=3,UART_ADDRESS_WIDTH=4) 
//

module \servo(DEV_ID=3,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_180, 
            n29239, n29762, n29196, C_5_c_c, n29225, n8720) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_180;
    input n29239;
    input n29762;
    input n29196;
    input C_5_c_c;
    input n29225;
    output n8720;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    FD1P3IX mode_60 (.D(n29762), .SP(clk_enable_180), .CD(n29239), .CK(clk), 
            .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=418, LSE_RLINE=453 */ ;   // c:/s_links/sources/slot_cards/servo.v(66[8] 74[4])
    defparam mode_60.GSR = "DISABLED";
    LUT4 i22817_3_lut_4_lut (.A(mode), .B(n29196), .C(C_5_c_c), .D(n29225), 
         .Z(n8720)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;   // c:/s_links/sources/slot_cards/servo.v(61[19:72])
    defparam i22817_3_lut_4_lut.init = 16'hfd00;
    
endmodule
//
// Verilog Description of module \servo(DEV_ID=1,UART_ADDRESS_WIDTH=4) 
//

module \servo(DEV_ID=1,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_184, 
            n29239, n29762, n29202, C_5_c_c, n29237, n8777) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_184;
    input n29239;
    input n29762;
    input n29202;
    input C_5_c_c;
    input n29237;
    output n8777;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    FD1P3IX mode_60 (.D(n29762), .SP(clk_enable_184), .CD(n29239), .CK(clk), 
            .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=418, LSE_RLINE=453 */ ;   // c:/s_links/sources/slot_cards/servo.v(66[8] 74[4])
    defparam mode_60.GSR = "DISABLED";
    LUT4 i22807_3_lut_4_lut (.A(mode), .B(n29202), .C(C_5_c_c), .D(n29237), 
         .Z(n8777)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;   // c:/s_links/sources/slot_cards/servo.v(61[19:72])
    defparam i22807_3_lut_4_lut.init = 16'hfd00;
    
endmodule
//
// Verilog Description of module \servo(DEV_ID=2,UART_ADDRESS_WIDTH=4) 
//

module \servo(DEV_ID=2,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_181, 
            n29239, n29762, n29194, C_5_c_c, n29233, n8749) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_181;
    input n29239;
    input n29762;
    input n29194;
    input C_5_c_c;
    input n29233;
    output n8749;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    FD1P3IX mode_60 (.D(n29762), .SP(clk_enable_181), .CD(n29239), .CK(clk), 
            .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=418, LSE_RLINE=453 */ ;   // c:/s_links/sources/slot_cards/servo.v(66[8] 74[4])
    defparam mode_60.GSR = "DISABLED";
    LUT4 i22812_3_lut_4_lut (.A(mode), .B(n29194), .C(C_5_c_c), .D(n29233), 
         .Z(n8749)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;   // c:/s_links/sources/slot_cards/servo.v(61[19:72])
    defparam i22812_3_lut_4_lut.init = 16'hfd00;
    
endmodule
//
// Verilog Description of module \servo(DEV_ID=5,UART_ADDRESS_WIDTH=4) 
//

module \servo(DEV_ID=5,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_175, 
            n29239, n29762, n29199, C_5_c_c, n29220, n8661) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_175;
    input n29239;
    input n29762;
    input n29199;
    input C_5_c_c;
    input n29220;
    output n8661;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    FD1P3IX mode_60 (.D(n29762), .SP(clk_enable_175), .CD(n29239), .CK(clk), 
            .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=418, LSE_RLINE=453 */ ;   // c:/s_links/sources/slot_cards/servo.v(66[8] 74[4])
    defparam mode_60.GSR = "DISABLED";
    LUT4 i22840_3_lut_4_lut (.A(mode), .B(n29199), .C(C_5_c_c), .D(n29220), 
         .Z(n8661)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;   // c:/s_links/sources/slot_cards/servo.v(61[19:72])
    defparam i22840_3_lut_4_lut.init = 16'hfd00;
    
endmodule
//
// Verilog Description of module \servo(UART_ADDRESS_WIDTH=4) 
//

module \servo(UART_ADDRESS_WIDTH=4)  (mode, n29160, C_5_c_c, n29260, 
            n8805, clk, clk_enable_186, n29239, n29762) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input n29160;
    input C_5_c_c;
    input n29260;
    output n8805;
    input clk;
    input clk_enable_186;
    input n29239;
    input n29762;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    LUT4 i22796_3_lut_4_lut (.A(mode), .B(n29160), .C(C_5_c_c), .D(n29260), 
         .Z(n8805)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;   // c:/s_links/sources/slot_cards/servo.v(61[19:72])
    defparam i22796_3_lut_4_lut.init = 16'hfd00;
    FD1P3IX mode_60 (.D(n29762), .SP(clk_enable_186), .CD(n29239), .CK(clk), 
            .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=418, LSE_RLINE=453 */ ;   // c:/s_links/sources/slot_cards/servo.v(66[8] 74[4])
    defparam mode_60.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \servo(DEV_ID=4,UART_ADDRESS_WIDTH=4) 
//

module \servo(DEV_ID=4,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_178, 
            n29239, n29762, n29204, C_5_c_c, n29224, n8689) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_178;
    input n29239;
    input n29762;
    input n29204;
    input C_5_c_c;
    input n29224;
    output n8689;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    FD1P3IX mode_60 (.D(n29762), .SP(clk_enable_178), .CD(n29239), .CK(clk), 
            .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=418, LSE_RLINE=453 */ ;   // c:/s_links/sources/slot_cards/servo.v(66[8] 74[4])
    defparam mode_60.GSR = "DISABLED";
    LUT4 i22835_3_lut_4_lut (.A(mode), .B(n29204), .C(C_5_c_c), .D(n29224), 
         .Z(n8689)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;   // c:/s_links/sources/slot_cards/servo.v(61[19:72])
    defparam i22835_3_lut_4_lut.init = 16'hfd00;
    
endmodule
//
// Verilog Description of module \otm_dac(DEV_ID=3) 
//

module \otm_dac(DEV_ID=3)  (NSL, n29317, mode, n8717, clk, clk_enable_193, 
            n29239, \spi_data_r[0] , clk_enable_204, n29214, n29127, 
            n27259, \spi_addr_r[1] , n29084, n29254, n27286, reset_r_N_4813, 
            n29162, n29085) /* synthesis syn_module_defined=1 */ ;
    input NSL;
    input n29317;
    output mode;
    output n8717;
    input clk;
    input clk_enable_193;
    input n29239;
    input \spi_data_r[0] ;
    input clk_enable_204;
    input n29214;
    input n29127;
    input n27259;
    input \spi_addr_r[1] ;
    output n29084;
    input n29254;
    input n27286;
    output reset_r_N_4813;
    input n29162;
    output n29085;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    wire LASER_CNTRL_r;
    
    LUT4 Select_3935_i7_4_lut (.A(NSL), .B(LASER_CNTRL_r), .C(n29317), 
         .D(mode), .Z(n8717)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam Select_3935_i7_4_lut.init = 16'heca0;
    FD1P3IX mode_30 (.D(\spi_data_r[0] ), .SP(clk_enable_193), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=577, LSE_RLINE=595 */ ;   // c:/s_links/sources/otm_dac.v(36[8] 44[4])
    defparam mode_30.GSR = "DISABLED";
    FD1P3IX LASER_CNTRL_r_31 (.D(\spi_data_r[0] ), .SP(clk_enable_204), 
            .CD(n29239), .CK(clk), .Q(LASER_CNTRL_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=577, LSE_RLINE=595 */ ;   // c:/s_links/sources/otm_dac.v(47[8] 55[4])
    defparam LASER_CNTRL_r_31.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_356_3_lut_4_lut (.A(n29214), .B(n29127), .C(n27259), 
         .D(\spi_addr_r[1] ), .Z(n29084)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_rep_356_3_lut_4_lut.init = 16'h0040;
    LUT4 i2_3_lut_4_lut (.A(n29214), .B(n29127), .C(n29254), .D(n27286), 
         .Z(reset_r_N_4813)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_rep_357_3_lut_4_lut (.A(n29214), .B(n29127), .C(n29162), 
         .D(\spi_addr_r[1] ), .Z(n29085)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_rep_357_3_lut_4_lut.init = 16'h0040;
    
endmodule
//
// Verilog Description of module \shutter(DEV_ID=1,UART_ADDRESS_WIDTH=4) 
//

module \shutter(DEV_ID=1,UART_ADDRESS_WIDTH=4)  (mode_adj_554, n29237, \quad_homing[1] , 
            n27636, n26963, n12716, pin_io_out_14, \pin_intrpt[5] , 
            pin_io_out_12, \pin_intrpt[3] , reset_r, n1, \cs_decoded[2] , 
            n2, n29198, pin_io_out_13, \pin_intrpt[4] , mode, clk, 
            clk_enable_179, n29239, \spi_data_r[0] , n8898) /* synthesis syn_module_defined=1 */ ;
    input [2:0]mode_adj_554;
    output n29237;
    input \quad_homing[1] ;
    input n27636;
    output n26963;
    output n12716;
    input pin_io_out_14;
    output \pin_intrpt[5] ;
    input pin_io_out_12;
    output \pin_intrpt[3] ;
    input reset_r;
    output n1;
    input \cs_decoded[2] ;
    output n2;
    output n29198;
    input pin_io_out_13;
    output \pin_intrpt[4] ;
    output mode;
    input clk;
    input clk_enable_179;
    input n29239;
    input \spi_data_r[0] ;
    output n8898;
    
    wire \pin_intrpt[5]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[5] */ ;   // c:/s_links/sources/mcm_top.v(102[46:56])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    LUT4 i22721_2_lut_rep_509 (.A(mode_adj_554[1]), .B(mode_adj_554[2]), 
         .Z(n29237)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i22721_2_lut_rep_509.init = 16'h1111;
    LUT4 i2_3_lut_4_lut (.A(mode_adj_554[1]), .B(mode_adj_554[2]), .C(\quad_homing[1] ), 
         .D(n27636), .Z(n26963)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;
    defparam i2_3_lut_4_lut.init = 16'hf1ff;
    LUT4 i3_3_lut_4_lut (.A(mode_adj_554[1]), .B(mode_adj_554[2]), .C(\quad_homing[1] ), 
         .D(n27636), .Z(n12716)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;
    defparam i3_3_lut_4_lut.init = 16'h0e00;
    LUT4 i4190_2_lut_3_lut (.A(mode_adj_554[1]), .B(mode_adj_554[2]), .C(pin_io_out_14), 
         .Z(\pin_intrpt[5] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i4190_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_4112_i1_2_lut_3_lut (.A(mode_adj_554[1]), .B(mode_adj_554[2]), 
         .C(pin_io_out_12), .Z(\pin_intrpt[3] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4112_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_4010_i1_2_lut_3_lut (.A(mode_adj_554[1]), .B(mode_adj_554[2]), 
         .C(reset_r), .Z(n1)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4010_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_3997_i2_2_lut_3_lut (.A(mode_adj_554[1]), .B(mode_adj_554[2]), 
         .C(\cs_decoded[2] ), .Z(n2)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_3997_i2_2_lut_3_lut.init = 16'he0e0;
    LUT4 i2_2_lut_rep_470_3_lut (.A(mode_adj_554[1]), .B(mode_adj_554[2]), 
         .C(mode_adj_554[0]), .Z(n29198)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_2_lut_rep_470_3_lut.init = 16'hfefe;
    LUT4 Select_4111_i1_2_lut_3_lut (.A(mode_adj_554[1]), .B(mode_adj_554[2]), 
         .C(pin_io_out_13), .Z(\pin_intrpt[4] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4111_i1_2_lut_3_lut.init = 16'he0e0;
    FD1P3IX mode_160 (.D(\spi_data_r[0] ), .SP(clk_enable_179), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=508, LSE_RLINE=540 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(81[8] 89[4])
    defparam mode_160.GSR = "DISABLED";
    LUT4 i4152_1_lut (.A(mode_adj_554[2]), .Z(n8898)) /* synthesis lut_function=(!(A)) */ ;
    defparam i4152_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module \peizo_elliptec(DEV_ID=7,UART_ADDRESS_WIDTH=4) 
//

module \peizo_elliptec(DEV_ID=7,UART_ADDRESS_WIDTH=4)  (clk, clk_enable_194, 
            n29239, \spi_data_r[0] , C_1_c_0, n29313, C_2_c_1, tx_N_6443) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input clk_enable_194;
    input n29239;
    input \spi_data_r[0] ;
    input C_1_c_0;
    input n29313;
    input C_2_c_1;
    output tx_N_6443;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    wire mode;
    
    FD1P3IX mode_26 (.D(\spi_data_r[0] ), .SP(clk_enable_194), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=602, LSE_RLINE=622 */ ;   // c:/s_links/sources/slot_cards/peizo_elliptec.v(36[8] 44[4])
    defparam mode_26.GSR = "DISABLED";
    LUT4 i22694_4_lut (.A(mode), .B(C_1_c_0), .C(n29313), .D(C_2_c_1), 
         .Z(tx_N_6443)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;   // c:/s_links/sources/slot_cards/peizo_elliptec.v(30[8:10])
    defparam i22694_4_lut.init = 16'hdfff;
    
endmodule
//
// Verilog Description of module \shutter(UART_ADDRESS_WIDTH=4) 
//

module \shutter(UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_189, n29239, 
            \spi_data_r[0] , \mode[1] , \mode[2] , n29260, \quad_homing[0] , 
            pin_io_out_4, n5, pin_io_out_2, \pin_intrpt[0] , reset_r, 
            n1, \cs_decoded[0] , n2, \mode[2]_derived_32 , pin_io_out_3, 
            \pin_intrpt[1] , n29160, mode_adj_553, n29201, n31, n27471, 
            n29089, n29254, n29083, resetn_c, clk_enable_198, n29214, 
            n29118, \spi_addr_r[1] , n27256, reset_r_N_4474, n19084, 
            \spi_cmd_r[1] , \spi_cmd_r[3] , n29082, n29182, \spi_cmd_r[0] , 
            n29130, n65, n27, \spi_addr_r[2] , n27283, clk_enable_164, 
            n29174, n29127, n27285, n29104, n29251, n29256, n29102, 
            n19233, n29100, n29096, n13074, clk_enable_173) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_189;
    input n29239;
    input \spi_data_r[0] ;
    input \mode[1] ;
    input \mode[2] ;
    output n29260;
    input \quad_homing[0] ;
    input pin_io_out_4;
    output n5;
    input pin_io_out_2;
    output \pin_intrpt[0] ;
    input reset_r;
    output n1;
    input \cs_decoded[0] ;
    output n2;
    output \mode[2]_derived_32 ;
    input pin_io_out_3;
    output \pin_intrpt[1] ;
    input n29160;
    input mode_adj_553;
    input n29201;
    input n31;
    output n27471;
    input n29089;
    input n29254;
    input n29083;
    input resetn_c;
    output clk_enable_198;
    input n29214;
    input n29118;
    input \spi_addr_r[1] ;
    input n27256;
    output reset_r_N_4474;
    input n19084;
    input \spi_cmd_r[1] ;
    input \spi_cmd_r[3] ;
    output n29082;
    input n29182;
    input \spi_cmd_r[0] ;
    input n29130;
    output n65;
    input n27;
    input \spi_addr_r[2] ;
    input n27283;
    output clk_enable_164;
    input n29174;
    input n29127;
    output n27285;
    output n29104;
    input n29251;
    input n29256;
    output n29102;
    input n19233;
    output n29100;
    input n29096;
    input n13074;
    output clk_enable_173;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire \mode[2]_derived_32  /* synthesis is_clock=1, SET_AS_NETWORK=\stepper_ins[0].u_stepper/mode[2]_derived_32 */ ;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    FD1P3IX mode_160 (.D(\spi_data_r[0] ), .SP(clk_enable_189), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=508, LSE_RLINE=540 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(81[8] 89[4])
    defparam mode_160.GSR = "DISABLED";
    LUT4 i22708_2_lut_rep_532 (.A(\mode[1] ), .B(\mode[2] ), .Z(n29260)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i22708_2_lut_rep_532.init = 16'h1111;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\mode[1] ), .B(\mode[2] ), .C(\quad_homing[0] ), 
         .D(pin_io_out_4), .Z(n5)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 Select_4114_i1_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(pin_io_out_2), 
         .Z(\pin_intrpt[0] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4114_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_4038_i1_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(reset_r), 
         .Z(n1)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4038_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_4025_i2_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(\cs_decoded[0] ), 
         .Z(n2)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4025_i2_2_lut_3_lut.init = 16'he0e0;
    LUT4 i4189_2_lut_rep_455_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(pin_io_out_4), 
         .Z(\mode[2]_derived_32 )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i4189_2_lut_rep_455_3_lut.init = 16'he0e0;
    LUT4 Select_4113_i1_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(pin_io_out_3), 
         .Z(\pin_intrpt[1] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4113_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 i1_4_lut (.A(n29160), .B(mode_adj_553), .C(n29201), .D(n31), 
         .Z(n27471)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(76[18:71])
    defparam i1_4_lut.init = 16'h5554;
    LUT4 i1_3_lut_4_lut (.A(n29089), .B(n29254), .C(n29083), .D(resetn_c), 
         .Z(clk_enable_198)) /* synthesis lut_function=(!(((C (D))+!B)+!A)) */ ;   // c:/s_links/sources/status_led.v(35[30:38])
    defparam i1_3_lut_4_lut.init = 16'h0888;
    LUT4 i2_3_lut_4_lut (.A(n29214), .B(n29118), .C(\spi_addr_r[1] ), 
         .D(n27256), .Z(reset_r_N_4474)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_rep_354_4_lut (.A(n19084), .B(\spi_cmd_r[1] ), .C(n29118), 
         .D(\spi_cmd_r[3] ), .Z(n29082)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_rep_354_4_lut.init = 16'h4000;
    LUT4 i3_4_lut (.A(\spi_addr_r[1] ), .B(n29182), .C(\spi_cmd_r[0] ), 
         .D(n29130), .Z(n65)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i3_4_lut.init = 16'h2000;
    LUT4 i3_4_lut_adj_969 (.A(n27), .B(\spi_addr_r[2] ), .C(n29118), .D(n27283), 
         .Z(clk_enable_164)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(35[30:38])
    defparam i3_4_lut_adj_969.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_970 (.A(n29174), .B(n29127), .C(n27283), 
         .D(n29214), .Z(n27285)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_970.init = 16'h0080;
    LUT4 i2_3_lut_rep_376_4_lut (.A(n29174), .B(n29127), .C(\spi_cmd_r[1] ), 
         .D(n19084), .Z(n29104)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_rep_376_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_374_4_lut (.A(\spi_cmd_r[0] ), .B(n29251), .C(n29130), 
         .D(n29256), .Z(n29102)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_374_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_372_4_lut (.A(\spi_cmd_r[0] ), .B(n29251), .C(n29130), 
         .D(n19233), .Z(n29100)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_372_4_lut.init = 16'h0010;
    LUT4 i4960_3_lut_4_lut (.A(\spi_cmd_r[3] ), .B(n29104), .C(n29096), 
         .D(n13074), .Z(clk_enable_173)) /* synthesis lut_function=(!(((C (D))+!B)+!A)) */ ;
    defparam i4960_3_lut_4_lut.init = 16'h0888;
    
endmodule
//
// Verilog Description of module \piezo(DEV_ID=1,UART_ADDRESS_WIDTH=4) 
//

module \piezo(DEV_ID=1,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_187, 
            n29239, \spi_data_r[0] , n29282, n29284, n29237, mode_adj_552, 
            OW_ID_N_4464, C_1_c_0, C_2_c_1, mode_adj_549, n29313, 
            n29158, mode_adj_550, n29157, n13, n27483, \cs_decoded[3] , 
            n2, n8908, digital_output_r, n26533, OW_ID_N_4462, C_5_c_c, 
            n29202, n13615, mode_adj_551, n29306, n29315, n8795) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_187;
    input n29239;
    input \spi_data_r[0] ;
    output n29282;
    input n29284;
    input n29237;
    input [2:0]mode_adj_552;
    output OW_ID_N_4464;
    input C_1_c_0;
    input C_2_c_1;
    input mode_adj_549;
    input n29313;
    output n29158;
    input mode_adj_550;
    output n29157;
    input n13;
    output n27483;
    input \cs_decoded[3] ;
    output n2;
    output n8908;
    input digital_output_r;
    output n26533;
    input OW_ID_N_4462;
    input C_5_c_c;
    input n29202;
    output n13615;
    input mode_adj_551;
    output n29306;
    input n29315;
    output n8795;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    FD1P3IX mode_38 (.D(\spi_data_r[0] ), .SP(clk_enable_187), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=632, LSE_RLINE=661 */ ;   // c:/s_links/sources/slot_cards/piezo.v(55[8] 63[4])
    defparam mode_38.GSR = "DISABLED";
    LUT4 OW_ID_I_125_2_lut_3_lut_4_lut (.A(n29282), .B(n29284), .C(n29237), 
         .D(mode_adj_552[0]), .Z(OW_ID_N_4464)) /* synthesis lut_function=(!(A+(B+!((D)+!C)))) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam OW_ID_I_125_2_lut_3_lut_4_lut.init = 16'h1101;
    LUT4 equal_272_i5_2_lut_rep_554 (.A(C_1_c_0), .B(C_2_c_1), .Z(n29282)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam equal_272_i5_2_lut_rep_554.init = 16'heeee;
    LUT4 OW_ID_I_275_2_lut_rep_430_3_lut_4_lut (.A(C_1_c_0), .B(C_2_c_1), 
         .C(mode_adj_549), .D(n29313), .Z(n29158)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam OW_ID_I_275_2_lut_rep_430_3_lut_4_lut.init = 16'h1000;
    LUT4 OW_ID_I_259_2_lut_rep_429_3_lut_4_lut (.A(C_1_c_0), .B(C_2_c_1), 
         .C(mode_adj_550), .D(n29284), .Z(n29157)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam OW_ID_I_259_2_lut_rep_429_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_3_lut_4_lut (.A(C_1_c_0), .B(C_2_c_1), .C(n13), .D(n29284), 
         .Z(n27483)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 Select_4007_i2_2_lut (.A(\cs_decoded[3] ), .B(mode), .Z(n2)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4007_i2_2_lut.init = 16'h8888;
    LUT4 i4157_1_lut (.A(mode), .Z(n8908)) /* synthesis lut_function=(!(A)) */ ;
    defparam i4157_1_lut.init = 16'h5555;
    LUT4 i3_4_lut (.A(mode_adj_552[2]), .B(mode_adj_552[0]), .C(digital_output_r), 
         .D(mode_adj_552[1]), .Z(n26533)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i3_4_lut.init = 16'h4000;
    LUT4 i22799_4_lut (.A(OW_ID_N_4462), .B(n13), .C(C_5_c_c), .D(n29202), 
         .Z(n13615)) /* synthesis lut_function=(!(A+!((C+(D))+!B))) */ ;
    defparam i22799_4_lut.init = 16'h5551;
    LUT4 i4014_2_lut_rep_578 (.A(mode_adj_551), .B(mode), .Z(n29306)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/piezo.v(46[8:14])
    defparam i4014_2_lut_rep_578.init = 16'heeee;
    LUT4 i22710_2_lut_2_lut_3_lut_4_lut (.A(mode_adj_551), .B(mode), .C(n29315), 
         .D(mode_adj_552[0]), .Z(n8795)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // c:/s_links/sources/slot_cards/piezo.v(46[8:14])
    defparam i22710_2_lut_2_lut_3_lut_4_lut.init = 16'h1011;
    
endmodule
//
// Verilog Description of module \piezo(UART_ADDRESS_WIDTH=4) 
//

module \piezo(UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_192, n29239, 
            \spi_data_r[0] , \spi_cmd_r[3] , n29251, \spi_addr_r[1] , 
            n29214, n29124, mode_adj_548, digital_output_r, n26535, 
            n26561, n27, \spi_addr_r[2] , n29161, n29169, n29216, 
            n27225, \spi_addr_r[0] , n19084, n29286, n29123, n29287, 
            n29101, \cs_decoded[1] , n2, n8922, C_5_c_c, n22, C_4_c_3, 
            n29200, n3, n29307, \spi_cmd_r[1] , n27240, mode_adj_547, 
            n29309, \spi_cmd_r[2] , n29288, n65, n27234) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_192;
    input n29239;
    input \spi_data_r[0] ;
    input \spi_cmd_r[3] ;
    input n29251;
    input \spi_addr_r[1] ;
    output n29214;
    output n29124;
    input [2:0]mode_adj_548;
    input digital_output_r;
    output n26535;
    output n26561;
    input n27;
    input \spi_addr_r[2] ;
    output n29161;
    output n29169;
    input n29216;
    output n27225;
    input \spi_addr_r[0] ;
    output n19084;
    output n29286;
    input n29123;
    input n29287;
    output n29101;
    input \cs_decoded[1] ;
    output n2;
    output n8922;
    input C_5_c_c;
    input n22;
    input C_4_c_3;
    input n29200;
    output n3;
    output n29307;
    input \spi_cmd_r[1] ;
    output n27240;
    input mode_adj_547;
    output n29309;
    input \spi_cmd_r[2] ;
    input n29288;
    output n65;
    output n27234;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    wire n26997;
    
    FD1P3IX mode_38 (.D(\spi_data_r[0] ), .SP(clk_enable_192), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=632, LSE_RLINE=661 */ ;   // c:/s_links/sources/slot_cards/piezo.v(55[8] 63[4])
    defparam mode_38.GSR = "DISABLED";
    LUT4 i14093_2_lut_rep_396_3_lut_4_lut (.A(\spi_cmd_r[3] ), .B(n29251), 
         .C(\spi_addr_r[1] ), .D(n29214), .Z(n29124)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14093_2_lut_rep_396_3_lut_4_lut.init = 16'hfffe;
    LUT4 i3_3_lut_4_lut (.A(mode_adj_548[0]), .B(mode_adj_548[1]), .C(digital_output_r), 
         .D(mode_adj_548[2]), .Z(n26535)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i3_3_lut_4_lut.init = 16'h0080;
    LUT4 i22794_3_lut_4_lut (.A(mode_adj_548[0]), .B(mode_adj_548[1]), .C(n26997), 
         .D(mode_adj_548[2]), .Z(n26561)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A (C))) */ ;
    defparam i22794_3_lut_4_lut.init = 16'h0f07;
    LUT4 i13886_2_lut_rep_486 (.A(n27), .B(\spi_addr_r[2] ), .Z(n29214)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13886_2_lut_rep_486.init = 16'heeee;
    LUT4 i1_2_lut_rep_433_3_lut (.A(n27), .B(\spi_addr_r[2] ), .C(\spi_addr_r[1] ), 
         .Z(n29161)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_433_3_lut.init = 16'h1010;
    LUT4 i14091_2_lut_rep_441_3_lut (.A(n27), .B(\spi_addr_r[2] ), .C(\spi_addr_r[1] ), 
         .Z(n29169)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i14091_2_lut_rep_441_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n27), .B(\spi_addr_r[2] ), .C(n29216), 
         .D(\spi_addr_r[1] ), .Z(n27225)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i14157_2_lut_3_lut_4_lut (.A(n27), .B(\spi_addr_r[2] ), .C(\spi_addr_r[0] ), 
         .D(\spi_addr_r[1] ), .Z(n19084)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14157_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i22424_2_lut_rep_558 (.A(\spi_addr_r[1] ), .B(\spi_cmd_r[3] ), 
         .Z(n29286)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22424_2_lut_rep_558.init = 16'heeee;
    LUT4 i2_3_lut_rep_373_4_lut (.A(\spi_addr_r[1] ), .B(\spi_cmd_r[3] ), 
         .C(n29123), .D(n29287), .Z(n29101)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_3_lut_rep_373_4_lut.init = 16'h1000;
    LUT4 Select_4035_i2_2_lut (.A(\cs_decoded[1] ), .B(mode), .Z(n2)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4035_i2_2_lut.init = 16'h8888;
    LUT4 i4164_1_lut (.A(mode), .Z(n8922)) /* synthesis lut_function=(!(A)) */ ;
    defparam i4164_1_lut.init = 16'h5555;
    LUT4 i3_4_lut (.A(C_5_c_c), .B(n22), .C(C_4_c_3), .D(n29200), .Z(n26997)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i3_4_lut.init = 16'h0400;
    LUT4 i1_1_lut (.A(mode_adj_548[2]), .Z(n3)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_rep_579 (.A(\spi_addr_r[1] ), .B(\spi_cmd_r[3] ), .Z(n29307)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/slot_cards/piezo.v(58[15:52])
    defparam i1_2_lut_rep_579.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_4_lut_adj_967 (.A(\spi_addr_r[1] ), .B(\spi_cmd_r[3] ), 
         .C(\spi_addr_r[0] ), .D(\spi_cmd_r[1] ), .Z(n27240)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/s_links/sources/slot_cards/piezo.v(58[15:52])
    defparam i1_2_lut_3_lut_4_lut_adj_967.init = 16'h0200;
    LUT4 i4042_2_lut_rep_581 (.A(mode_adj_547), .B(mode), .Z(n29309)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/piezo.v(46[8:14])
    defparam i4042_2_lut_rep_581.init = 16'heeee;
    LUT4 i3_4_lut_adj_968 (.A(\spi_cmd_r[2] ), .B(n29123), .C(n29288), 
         .D(n65), .Z(n27234)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i3_4_lut_adj_968.init = 16'h4000;
    LUT4 i1_2_lut (.A(\spi_addr_r[1] ), .B(\spi_cmd_r[3] ), .Z(n65)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    
endmodule
//
// Verilog Description of module \piezo(DEV_ID=2,UART_ADDRESS_WIDTH=4) 
//

module \piezo(DEV_ID=2,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_185, 
            n29239, n29762, \cs_decoded[5] , n2, n8894, mode_adj_546, 
            digital_output_r, n26531, n26549, n27590, C_2_c_1, C_1_c_0, 
            n22, n8884) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_185;
    input n29239;
    input n29762;
    input \cs_decoded[5] ;
    output n2;
    output n8894;
    input [2:0]mode_adj_546;
    input digital_output_r;
    output n26531;
    output n26549;
    input n27590;
    input C_2_c_1;
    input C_1_c_0;
    input n22;
    output n8884;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    wire n27263;
    
    FD1P3IX mode_38 (.D(n29762), .SP(clk_enable_185), .CD(n29239), .CK(clk), 
            .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=632, LSE_RLINE=661 */ ;   // c:/s_links/sources/slot_cards/piezo.v(55[8] 63[4])
    defparam mode_38.GSR = "DISABLED";
    LUT4 Select_3979_i2_2_lut (.A(\cs_decoded[5] ), .B(mode), .Z(n2)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_3979_i2_2_lut.init = 16'h8888;
    LUT4 i4150_1_lut (.A(mode), .Z(n8894)) /* synthesis lut_function=(!(A)) */ ;
    defparam i4150_1_lut.init = 16'h5555;
    LUT4 i3_4_lut (.A(mode_adj_546[2]), .B(mode_adj_546[0]), .C(digital_output_r), 
         .D(mode_adj_546[1]), .Z(n26531)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i3_4_lut.init = 16'h4000;
    LUT4 i22810_4_lut (.A(mode_adj_546[1]), .B(n27263), .C(mode_adj_546[2]), 
         .D(mode_adj_546[0]), .Z(n26549)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B))) */ ;
    defparam i22810_4_lut.init = 16'h3133;
    LUT4 i2_4_lut (.A(n27590), .B(C_2_c_1), .C(C_1_c_0), .D(n22), .Z(n27263)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_4_lut.init = 16'h1000;
    LUT4 i1_1_lut (.A(mode_adj_546[2]), .Z(n8884)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module \piezo(DEV_ID=3,UART_ADDRESS_WIDTH=4) 
//

module \piezo(DEV_ID=3,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_183, 
            n29239, n29762, n29203, n29300, mode_adj_544, pin_io_out_35, 
            n26972, \cs_decoded[7] , n2, n8880, mode_adj_545, digital_output_r, 
            n26529, n26565, n27590, C_1_c_0, C_2_c_1, n29149, n8870) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_183;
    input n29239;
    input n29762;
    input n29203;
    input n29300;
    input mode_adj_544;
    input pin_io_out_35;
    output n26972;
    input \cs_decoded[7] ;
    output n2;
    output n8880;
    input [2:0]mode_adj_545;
    input digital_output_r;
    output n26529;
    output n26565;
    input n27590;
    input C_1_c_0;
    input C_2_c_1;
    input n29149;
    output n8870;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    wire n27264;
    
    FD1P3IX mode_38 (.D(n29762), .SP(clk_enable_183), .CD(n29239), .CK(clk), 
            .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=632, LSE_RLINE=661 */ ;   // c:/s_links/sources/slot_cards/piezo.v(55[8] 63[4])
    defparam mode_38.GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut (.A(n29203), .B(n29300), .C(mode_adj_544), .D(pin_io_out_35), 
         .Z(n26972)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hfe00;
    LUT4 Select_3950_i2_2_lut (.A(\cs_decoded[7] ), .B(mode), .Z(n2)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_3950_i2_2_lut.init = 16'h8888;
    LUT4 i4143_1_lut (.A(mode), .Z(n8880)) /* synthesis lut_function=(!(A)) */ ;
    defparam i4143_1_lut.init = 16'h5555;
    LUT4 i3_4_lut (.A(mode_adj_545[2]), .B(mode_adj_545[0]), .C(digital_output_r), 
         .D(mode_adj_545[1]), .Z(n26529)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i3_4_lut.init = 16'h4000;
    LUT4 i22815_4_lut (.A(mode_adj_545[1]), .B(n27264), .C(mode_adj_545[2]), 
         .D(mode_adj_545[0]), .Z(n26565)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B))) */ ;
    defparam i22815_4_lut.init = 16'h3133;
    LUT4 i2_4_lut (.A(n27590), .B(C_1_c_0), .C(C_2_c_1), .D(n29149), 
         .Z(n27264)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_4_lut.init = 16'h1000;
    LUT4 i1_1_lut (.A(mode_adj_545[2]), .Z(n8870)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module \piezo(DEV_ID=4,UART_ADDRESS_WIDTH=4) 
//

module \piezo(DEV_ID=4,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_177, 
            n29239, n29762, mode_adj_543, digital_output_r, n26525, 
            C_4_c_3, n29200, pin_io_out_6, mode_adj_539, n7, C_3_c_2, 
            n29132, C_1_c_0, C_2_c_1, n29160, mode_adj_540, n29284, 
            n29150, n29196, n29202, n29204, C_5_c_c, n27590, n29194, 
            OW_ID_N_5482, mode_adj_541, n27189, mode_adj_542, \cs_decoded[9] , 
            n2, n8864, n26569, n8854) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_177;
    input n29239;
    input n29762;
    input [2:0]mode_adj_543;
    input digital_output_r;
    output n26525;
    input C_4_c_3;
    output n29200;
    input pin_io_out_6;
    input mode_adj_539;
    output n7;
    input C_3_c_2;
    output n29132;
    input C_1_c_0;
    input C_2_c_1;
    output n29160;
    input mode_adj_540;
    output n29284;
    output n29150;
    output n29196;
    output n29202;
    output n29204;
    input C_5_c_c;
    output n27590;
    output n29194;
    input OW_ID_N_5482;
    input mode_adj_541;
    output n27189;
    input mode_adj_542;
    input \cs_decoded[9] ;
    output n2;
    output n8864;
    output n26569;
    output n8854;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    wire n29264, n29283, n6;
    
    FD1P3IX mode_38 (.D(n29762), .SP(clk_enable_177), .CD(n29239), .CK(clk), 
            .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=632, LSE_RLINE=661 */ ;   // c:/s_links/sources/slot_cards/piezo.v(55[8] 63[4])
    defparam mode_38.GSR = "DISABLED";
    LUT4 i2_2_lut_rep_536 (.A(mode_adj_543[0]), .B(mode_adj_543[1]), .Z(n29264)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_rep_536.init = 16'h8888;
    LUT4 i3_3_lut_4_lut (.A(mode_adj_543[0]), .B(mode_adj_543[1]), .C(digital_output_r), 
         .D(mode_adj_543[2]), .Z(n26525)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i3_3_lut_4_lut.init = 16'h0080;
    LUT4 Select_3812_i7_2_lut_3_lut_4_lut (.A(C_4_c_3), .B(n29200), .C(pin_io_out_6), 
         .D(mode_adj_539), .Z(n7)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam Select_3812_i7_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 OW_ID_I_255_2_lut_rep_404_3_lut_4_lut (.A(n29283), .B(C_3_c_2), 
         .C(mode_adj_539), .D(C_4_c_3), .Z(n29132)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam OW_ID_I_255_2_lut_rep_404_3_lut_4_lut.init = 16'h0080;
    LUT4 i13603_2_lut_rep_555 (.A(C_1_c_0), .B(C_2_c_1), .Z(n29283)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13603_2_lut_rep_555.init = 16'h8888;
    LUT4 i22432_2_lut_rep_472_3_lut (.A(C_1_c_0), .B(C_2_c_1), .C(C_3_c_2), 
         .Z(n29200)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i22432_2_lut_rep_472_3_lut.init = 16'h8080;
    LUT4 i2_2_lut_rep_432_3_lut_4_lut (.A(C_1_c_0), .B(C_2_c_1), .C(C_4_c_3), 
         .D(C_3_c_2), .Z(n29160)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i2_2_lut_rep_432_3_lut_4_lut.init = 16'hf7ff;
    LUT4 OW_ID_I_271_2_lut_rep_422_3_lut_4_lut (.A(C_1_c_0), .B(C_2_c_1), 
         .C(mode_adj_540), .D(n29284), .Z(n29150)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam OW_ID_I_271_2_lut_rep_422_3_lut_4_lut.init = 16'h0080;
    LUT4 equal_284_i6_2_lut_rep_556 (.A(C_3_c_2), .B(C_4_c_3), .Z(n29284)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam equal_284_i6_2_lut_rep_556.init = 16'hbbbb;
    LUT4 i2_3_lut_rep_468_4_lut (.A(C_3_c_2), .B(C_4_c_3), .C(C_1_c_0), 
         .D(C_2_c_1), .Z(n29196)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam i2_3_lut_rep_468_4_lut.init = 16'hfbff;
    LUT4 equal_272_i7_2_lut_rep_474_3_lut_4_lut (.A(C_3_c_2), .B(C_4_c_3), 
         .C(C_2_c_1), .D(C_1_c_0), .Z(n29202)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam equal_272_i7_2_lut_rep_474_3_lut_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut_rep_476_3_lut_4_lut (.A(C_3_c_2), .B(C_4_c_3), .C(C_2_c_1), 
         .D(C_1_c_0), .Z(n29204)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam i1_2_lut_rep_476_3_lut_4_lut.init = 16'hbfff;
    LUT4 i22422_2_lut_3_lut (.A(C_3_c_2), .B(C_4_c_3), .C(C_5_c_c), .Z(n27590)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam i22422_2_lut_3_lut.init = 16'hfbfb;
    LUT4 i1_2_lut_rep_466_3_lut_4_lut (.A(C_3_c_2), .B(C_4_c_3), .C(C_1_c_0), 
         .D(C_2_c_1), .Z(n29194)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam i1_2_lut_rep_466_3_lut_4_lut.init = 16'hffbf;
    LUT4 i1_4_lut (.A(n29204), .B(OW_ID_N_5482), .C(n6), .D(mode_adj_541), 
         .Z(n27189)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;
    defparam i1_4_lut.init = 16'h5554;
    LUT4 i2_2_lut (.A(mode_adj_542), .B(mode), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 Select_3919_i2_2_lut (.A(\cs_decoded[9] ), .B(mode), .Z(n2)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_3919_i2_2_lut.init = 16'h8888;
    LUT4 i4135_1_lut (.A(mode), .Z(n8864)) /* synthesis lut_function=(!(A)) */ ;
    defparam i4135_1_lut.init = 16'h5555;
    LUT4 i22833_4_lut (.A(mode_adj_543[2]), .B(C_5_c_c), .C(n29264), .D(n27189), 
         .Z(n26569)) /* synthesis lut_function=(A (B+!(D))+!A !(B (C)+!B (C+(D)))) */ ;
    defparam i22833_4_lut.init = 16'h8caf;
    LUT4 i1_1_lut (.A(mode_adj_543[2]), .Z(n8854)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module \intrpt_ctrl(DEV_ID=5) 
//

module \intrpt_ctrl(DEV_ID=5)  (\spi_data_out_r_39__N_2927[0] , clk, \pin_intrpt[15] , 
            n29239, clear_intrpt, clear_intrpt_N_2994, intrpt_out_c_5, 
            intrpt_out_N_2990, n29757, \spi_data_out_r_39__N_2927[2] , 
            \mode[2]_derived_32 , \spi_data_out_r_39__N_2927[1] , \pin_intrpt[16] ) /* synthesis syn_module_defined=1 */ ;
    output \spi_data_out_r_39__N_2927[0] ;
    input clk;
    input \pin_intrpt[15] ;
    input n29239;
    output clear_intrpt;
    input clear_intrpt_N_2994;
    output intrpt_out_c_5;
    input intrpt_out_N_2990;
    input n29757;
    output \spi_data_out_r_39__N_2927[2] ;
    input \mode[2]_derived_32 ;
    output \spi_data_out_r_39__N_2927[1] ;
    input \pin_intrpt[16] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire \mode[2]_derived_32  /* synthesis is_clock=1, SET_AS_NETWORK=\stepper_ins[5].u_stepper/mode[2]_derived_32 */ ;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    wire [2:0]intrpt_in_reg;   // c:/s_links/sources/intrpt_ctrl.v(38[35:48])
    wire [2:0]intrpt_in_dly;   // c:/s_links/sources/intrpt_ctrl.v(39[36:49])
    
    wire assert_intrpt, intrpt_all_edges, n4;
    
    FD1S3AX spi_data_out_r_i1 (.D(\pin_intrpt[15] ), .CK(clk), .Q(\spi_data_out_r_39__N_2927[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i0 (.D(\pin_intrpt[15] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i0.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i0 (.D(intrpt_in_reg[0]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i0.GSR = "DISABLED";
    FD1S3IX clear_intrpt_317 (.D(clear_intrpt_N_2994), .CK(clk), .CD(n29239), 
            .Q(clear_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam clear_intrpt_317.GSR = "DISABLED";
    FD1S3IX assert_intrpt_316 (.D(intrpt_all_edges), .CK(clk), .CD(n29239), 
            .Q(assert_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(63[8] 73[4])
    defparam assert_intrpt_316.GSR = "DISABLED";
    FD1P3IX intrpt_out_359 (.D(n29757), .SP(assert_intrpt), .CD(intrpt_out_N_2990), 
            .CK(clk), .Q(intrpt_out_c_5)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(92[8] 99[4])
    defparam intrpt_out_359.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\mode[2]_derived_32 ), .CK(clk), .Q(\spi_data_out_r_39__N_2927[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\pin_intrpt[16] ), .CK(clk), .Q(\spi_data_out_r_39__N_2927[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i1 (.D(\pin_intrpt[16] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i2 (.D(\mode[2]_derived_32 ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i1 (.D(intrpt_in_reg[1]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i2 (.D(intrpt_in_reg[2]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i2.GSR = "DISABLED";
    LUT4 i2_3_lut (.A(intrpt_in_dly[0]), .B(n4), .C(intrpt_in_reg[0]), 
         .Z(intrpt_all_edges)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i2_3_lut.init = 16'hdede;
    LUT4 i1_4_lut (.A(intrpt_in_dly[1]), .B(intrpt_in_dly[2]), .C(intrpt_in_reg[1]), 
         .D(intrpt_in_reg[2]), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i1_4_lut.init = 16'h7bde;
    
endmodule
//
// Verilog Description of module \shutter(DEV_ID=6,UART_ADDRESS_WIDTH=4) 
//

module \shutter(DEV_ID=6,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_32, 
            n29239, \spi_data_r[0] , mode_adj_538, n29267, pin_io_out_64, 
            \pin_intrpt[20] , pin_io_out_62, \pin_intrpt[18] , pin_io_out_63, 
            \pin_intrpt[19] , reset_r, n1, \cs_decoded[12] , n2, n29190, 
            n8826) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_32;
    input n29239;
    input \spi_data_r[0] ;
    input [2:0]mode_adj_538;
    output n29267;
    input pin_io_out_64;
    output \pin_intrpt[20] ;
    input pin_io_out_62;
    output \pin_intrpt[18] ;
    input pin_io_out_63;
    output \pin_intrpt[19] ;
    input reset_r;
    output n1;
    input \cs_decoded[12] ;
    output n2;
    output n29190;
    output n8826;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire \pin_intrpt[20]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[20] */ ;   // c:/s_links/sources/mcm_top.v(102[46:56])
    
    FD1P3IX mode_160 (.D(\spi_data_r[0] ), .SP(clk_enable_32), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=508, LSE_RLINE=540 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(81[8] 89[4])
    defparam mode_160.GSR = "DISABLED";
    LUT4 i22788_2_lut_rep_539 (.A(mode_adj_538[1]), .B(mode_adj_538[2]), 
         .Z(n29267)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i22788_2_lut_rep_539.init = 16'h1111;
    LUT4 i4195_2_lut_3_lut (.A(mode_adj_538[1]), .B(mode_adj_538[2]), .C(pin_io_out_64), 
         .Z(\pin_intrpt[20] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i4195_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_4102_i1_2_lut_3_lut (.A(mode_adj_538[1]), .B(mode_adj_538[2]), 
         .C(pin_io_out_62), .Z(\pin_intrpt[18] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4102_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_4101_i1_2_lut_3_lut (.A(mode_adj_538[1]), .B(mode_adj_538[2]), 
         .C(pin_io_out_63), .Z(\pin_intrpt[19] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4101_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_3866_i1_2_lut_3_lut (.A(mode_adj_538[1]), .B(mode_adj_538[2]), 
         .C(reset_r), .Z(n1)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_3866_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_3853_i2_2_lut_3_lut (.A(mode_adj_538[1]), .B(mode_adj_538[2]), 
         .C(\cs_decoded[12] ), .Z(n2)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_3853_i2_2_lut_3_lut.init = 16'he0e0;
    LUT4 i2_2_lut_rep_462_3_lut (.A(mode_adj_538[1]), .B(mode_adj_538[2]), 
         .C(mode_adj_538[0]), .Z(n29190)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_2_lut_rep_462_3_lut.init = 16'hfefe;
    LUT4 i4116_1_lut (.A(mode_adj_538[2]), .Z(n8826)) /* synthesis lut_function=(!(A)) */ ;
    defparam i4116_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module \shutter(DEV_ID=5,UART_ADDRESS_WIDTH=4) 
//

module \shutter(DEV_ID=5,UART_ADDRESS_WIDTH=4)  (\mode[1] , \mode[2] , n29220, 
            \quad_homing[0] , pin_io_out_54, n27657, pin_io_out_52, 
            \pin_intrpt[15] , reset_r, n1, \cs_decoded[10] , n2, \mode[2]_derived_32 , 
            pin_io_out_53, \pin_intrpt[16] , mode, clk, clk_enable_172, 
            n29239, \spi_data_r[0] ) /* synthesis syn_module_defined=1 */ ;
    input \mode[1] ;
    input \mode[2] ;
    output n29220;
    input \quad_homing[0] ;
    input pin_io_out_54;
    output n27657;
    input pin_io_out_52;
    output \pin_intrpt[15] ;
    input reset_r;
    output n1;
    input \cs_decoded[10] ;
    output n2;
    output \mode[2]_derived_32 ;
    input pin_io_out_53;
    output \pin_intrpt[16] ;
    output mode;
    input clk;
    input clk_enable_172;
    input n29239;
    input \spi_data_r[0] ;
    
    wire \mode[2]_derived_32  /* synthesis is_clock=1, SET_AS_NETWORK=\stepper_ins[5].u_stepper/mode[2]_derived_32 */ ;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    LUT4 i22768_2_lut_rep_492 (.A(\mode[1] ), .B(\mode[2] ), .Z(n29220)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i22768_2_lut_rep_492.init = 16'h1111;
    LUT4 i22485_2_lut_3_lut_4_lut (.A(\mode[1] ), .B(\mode[2] ), .C(\quad_homing[0] ), 
         .D(pin_io_out_54), .Z(n27657)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i22485_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 Select_4104_i1_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(pin_io_out_52), 
         .Z(\pin_intrpt[15] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4104_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_3894_i1_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(reset_r), 
         .Z(n1)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_3894_i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 Select_3881_i2_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(\cs_decoded[10] ), 
         .Z(n2)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_3881_i2_2_lut_3_lut.init = 16'he0e0;
    LUT4 i4194_2_lut_rep_443_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(pin_io_out_54), 
         .Z(\mode[2]_derived_32 )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i4194_2_lut_rep_443_3_lut.init = 16'he0e0;
    LUT4 Select_4103_i1_2_lut_3_lut (.A(\mode[1] ), .B(\mode[2] ), .C(pin_io_out_53), 
         .Z(\pin_intrpt[16] )) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_4103_i1_2_lut_3_lut.init = 16'he0e0;
    FD1P3IX mode_160 (.D(\spi_data_r[0] ), .SP(clk_enable_172), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=508, LSE_RLINE=540 */ ;   // c:/s_links/sources/slot_cards/shutter_4.v(81[8] 89[4])
    defparam mode_160.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \io(DEV_ID=6,UART_ADDRESS_WIDTH=4) 
//

module \io(DEV_ID=6,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_191, 
            n29239, \spi_data_r[0] ) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_191;
    input n29239;
    input \spi_data_r[0] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    FD1P3IX mode_90 (.D(\spi_data_r[0] ), .SP(clk_enable_191), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=464, LSE_RLINE=496 */ ;   // c:/s_links/sources/slot_cards/slider_io.v(80[8] 88[4])
    defparam mode_90.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \status_led(DEV_ID=9) 
//

module \status_led(DEV_ID=9)  (clk, resetn_c, clk_enable_303, n29239, 
            \spi_data_r[0] , GND_net, \spi_data_out_r_39__N_770[0] , spi_data_out_r_39__N_810, 
            EM_STOP, led_sw_c, \spi_cmd_r[8] , n13265, \spi_cmd_r[14] , 
            \spi_cmd_r[11] , \spi_cmd_r[9] , \spi_cmd_r[13] , \spi_cmd_r[7] , 
            \spi_cmd_r[10] , spi_data_valid_r, \spi_cmd_r[12] , \spi_cmd_r[6] , 
            \spi_cmd_r[15] , \spi_data_r[11] , \spi_data_r[10] , \spi_data_r[9] , 
            \spi_data_r[8] , \spi_data_r[7] , \spi_data_r[6] , \spi_data_r[5] , 
            \spi_data_r[4] , \spi_data_r[3] , \spi_data_r[2] , \spi_data_r[1] , 
            n6, \spi_addr[3] , n27465, \spi_cmd[1] , \spi_addr[0] , 
            n13489, n26928) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input resetn_c;
    input clk_enable_303;
    input n29239;
    input \spi_data_r[0] ;
    input GND_net;
    output \spi_data_out_r_39__N_770[0] ;
    output spi_data_out_r_39__N_810;
    output EM_STOP;
    output led_sw_c;
    input \spi_cmd_r[8] ;
    output n13265;
    input \spi_cmd_r[14] ;
    input \spi_cmd_r[11] ;
    input \spi_cmd_r[9] ;
    input \spi_cmd_r[13] ;
    input \spi_cmd_r[7] ;
    input \spi_cmd_r[10] ;
    input spi_data_valid_r;
    input \spi_cmd_r[12] ;
    input \spi_cmd_r[6] ;
    input \spi_cmd_r[15] ;
    input \spi_data_r[11] ;
    input \spi_data_r[10] ;
    input \spi_data_r[9] ;
    input \spi_data_r[8] ;
    input \spi_data_r[7] ;
    input \spi_data_r[6] ;
    input \spi_data_r[5] ;
    input \spi_data_r[4] ;
    input \spi_data_r[3] ;
    input \spi_data_r[2] ;
    input \spi_data_r[1] ;
    input n6;
    input \spi_addr[3] ;
    input n27465;
    input \spi_cmd[1] ;
    input \spi_addr[0] ;
    input n13489;
    input n26928;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire [11:0]pwm_freq_cntr;   // c:/s_links/sources/status_led.v(36[30:43])
    
    wire n14284;
    wire [11:0]n53;
    wire [11:0]pwm_duty;   // c:/s_links/sources/status_led.v(35[30:38])
    
    wire n24970;
    wire [12:0]status_cntr;   // c:/s_links/sources/status_led.v(37[32:43])
    wire [12:0]n827;
    
    wire n24971, em_stop_flag, n13490, n29249, n14175, clk_enable_308, 
        n14229, n19611;
    wire [12:0]n141;
    
    wire n14283, n19475, pwm_out_N_893, clk_enable_205, n27015, n15, 
        n14, n29755, n27649, n27659, n18, n27614, n24972, n24968, 
        n24935, pwm_N_898, n24932;
    wire [12:0]pwm_N_899;
    
    wire n24933, n24934, n25205, n24969, n24973, n25204, n25203, 
        n25202, n25201, n25200, clk_enable_517, n25050, n25049, 
        n17, n22, n18_adj_7606, pwm_N_896, n25048, n25047, n20, 
        n14_adj_7607, n25046, n25045, n29219, n26939, n10, pwm, 
        n14160, n12, n14161, n4, n25288;
    
    FD1P3IX pwm_freq_cntr_2503__i1 (.D(n53[1]), .SP(resetn_c), .CD(n14284), 
            .CK(clk), .Q(pwm_freq_cntr[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503__i1.GSR = "DISABLED";
    FD1P3IX pwm_duty__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_303), .CD(n29239), 
            .CK(clk), .Q(pwm_duty[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i0.GSR = "DISABLED";
    CCU2D add_395_7 (.A0(status_cntr[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(status_cntr[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24970), .COUT(n24971), .S0(n827[5]), .S1(n827[6]));   // c:/s_links/sources/status_led.v(59[19:34])
    defparam add_395_7.INIT0 = 16'h5aaa;
    defparam add_395_7.INIT1 = 16'h5aaa;
    defparam add_395_7.INJECT1_0 = "NO";
    defparam add_395_7.INJECT1_1 = "NO";
    FD1S3AX spi_data_out_r_i1 (.D(em_stop_flag), .CK(clk), .Q(\spi_data_out_r_39__N_770[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(97[8] 111[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3IX i60_343 (.D(n29249), .CK(clk), .CD(n13490), .Q(spi_data_out_r_39__N_810)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(97[8] 111[4])
    defparam i60_343.GSR = "DISABLED";
    FD1S3AX em_stop_flag_383 (.D(n14175), .CK(clk), .Q(em_stop_flag)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(97[8] 111[4])
    defparam em_stop_flag_383.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_2503__i0 (.D(n53[0]), .SP(resetn_c), .CD(n14284), 
            .CK(clk), .Q(pwm_freq_cntr[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503__i0.GSR = "DISABLED";
    FD1P3IX status_cntr_i0_i1 (.D(n827[1]), .SP(clk_enable_308), .CD(n14229), 
            .CK(clk), .Q(status_cntr[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i1.GSR = "DISABLED";
    FD1P3IX status_cntr_i0_i2 (.D(n827[2]), .SP(clk_enable_308), .CD(n14229), 
            .CK(clk), .Q(status_cntr[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i2.GSR = "DISABLED";
    FD1P3IX status_cntr_i0_i3 (.D(n827[3]), .SP(clk_enable_308), .CD(n14229), 
            .CK(clk), .Q(status_cntr[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i3.GSR = "DISABLED";
    FD1P3JX status_cntr_i0_i4 (.D(n141[4]), .SP(clk_enable_308), .PD(n19611), 
            .CK(clk), .Q(status_cntr[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i4.GSR = "DISABLED";
    FD1P3IX status_cntr_i0_i5 (.D(n827[5]), .SP(clk_enable_308), .CD(n14229), 
            .CK(clk), .Q(status_cntr[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i5.GSR = "DISABLED";
    FD1P3JX status_cntr_i0_i6 (.D(n141[6]), .SP(clk_enable_308), .PD(n19611), 
            .CK(clk), .Q(status_cntr[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i6.GSR = "DISABLED";
    FD1P3JX status_cntr_i0_i7 (.D(n141[7]), .SP(clk_enable_308), .PD(n19611), 
            .CK(clk), .Q(status_cntr[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i7.GSR = "DISABLED";
    FD1P3JX status_cntr_i0_i8 (.D(n141[8]), .SP(clk_enable_308), .PD(n19611), 
            .CK(clk), .Q(status_cntr[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i8.GSR = "DISABLED";
    FD1P3JX status_cntr_i0_i9 (.D(n141[9]), .SP(clk_enable_308), .PD(n19611), 
            .CK(clk), .Q(status_cntr[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i9.GSR = "DISABLED";
    FD1P3JX status_cntr_i0_i10 (.D(n141[10]), .SP(clk_enable_308), .PD(n19611), 
            .CK(clk), .Q(status_cntr[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i10.GSR = "DISABLED";
    FD1P3IX status_cntr_i0_i11 (.D(n827[11]), .SP(clk_enable_308), .CD(n14229), 
            .CK(clk), .Q(status_cntr[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i11.GSR = "DISABLED";
    FD1P3IX status_cntr_i0_i12 (.D(n827[12]), .SP(clk_enable_308), .CD(n14229), 
            .CK(clk), .Q(status_cntr[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i12.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(n14283), .B(n827[4]), .Z(n141[4])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i22583_2_lut_rep_521 (.A(resetn_c), .B(EM_STOP), .Z(n29249)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/status_led.v(102[11] 110[5])
    defparam i22583_2_lut_rep_521.init = 16'h2222;
    LUT4 i9219_3_lut_4_lut (.A(resetn_c), .B(EM_STOP), .C(em_stop_flag), 
         .D(n13490), .Z(n14175)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(102[11] 110[5])
    defparam i9219_3_lut_4_lut.init = 16'hfddd;
    LUT4 i22896_2_lut_3_lut_4_lut (.A(n19475), .B(status_cntr[12]), .C(clk_enable_308), 
         .D(n14283), .Z(n14229)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam i22896_2_lut_3_lut_4_lut.init = 16'h80f0;
    LUT4 i9382_2_lut (.A(resetn_c), .B(n14283), .Z(n14284)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam i9382_2_lut.init = 16'h8888;
    FD1S3IX EM_STOP_338 (.D(pwm_out_N_893), .CK(clk), .CD(n29239), .Q(EM_STOP)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam EM_STOP_338.GSR = "DISABLED";
    FD1P3AX pwm_out_337 (.D(n27015), .SP(clk_enable_205), .CK(clk), .Q(led_sw_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_out_337.GSR = "DISABLED";
    LUT4 i8_4_lut (.A(n15), .B(pwm_freq_cntr[6]), .C(n14), .D(pwm_freq_cntr[1]), 
         .Z(n14283)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i8_4_lut.init = 16'h8000;
    LUT4 i6_4_lut (.A(pwm_freq_cntr[10]), .B(pwm_freq_cntr[8]), .C(pwm_freq_cntr[9]), 
         .D(pwm_freq_cntr[3]), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i6_4_lut.init = 16'h8000;
    LUT4 i14616_2_lut_rep_592 (.A(n19475), .B(status_cntr[12]), .Z(n29755)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14616_2_lut_rep_592.init = 16'h8888;
    LUT4 i14670_2_lut_2_lut_3_lut (.A(n19475), .B(status_cntr[12]), .C(resetn_c), 
         .Z(n19611)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i14670_2_lut_2_lut_3_lut.init = 16'h8080;
    LUT4 i5_3_lut (.A(n27649), .B(pwm_freq_cntr[5]), .C(pwm_freq_cntr[0]), 
         .Z(n14)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i5_3_lut.init = 16'h4040;
    LUT4 i22477_4_lut (.A(pwm_freq_cntr[4]), .B(pwm_freq_cntr[2]), .C(pwm_freq_cntr[7]), 
         .D(pwm_freq_cntr[11]), .Z(n27649)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22477_4_lut.init = 16'hfffe;
    LUT4 i10_4_lut (.A(n27659), .B(\spi_cmd_r[8] ), .C(n18), .D(n27614), 
         .Z(n13265)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i10_4_lut.init = 16'h0010;
    LUT4 i22487_4_lut (.A(\spi_cmd_r[14] ), .B(\spi_cmd_r[11] ), .C(\spi_cmd_r[9] ), 
         .D(\spi_cmd_r[13] ), .Z(n27659)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22487_4_lut.init = 16'hfffe;
    CCU2D add_395_9 (.A0(status_cntr[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(status_cntr[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24971), .COUT(n24972), .S0(n827[7]), .S1(n827[8]));   // c:/s_links/sources/status_led.v(59[19:34])
    defparam add_395_9.INIT0 = 16'h5aaa;
    defparam add_395_9.INIT1 = 16'h5aaa;
    defparam add_395_9.INJECT1_0 = "NO";
    defparam add_395_9.INJECT1_1 = "NO";
    CCU2D add_395_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(status_cntr[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24968), .S1(n827[0]));   // c:/s_links/sources/status_led.v(59[19:34])
    defparam add_395_1.INIT0 = 16'hF000;
    defparam add_395_1.INIT1 = 16'h5555;
    defparam add_395_1.INJECT1_0 = "NO";
    defparam add_395_1.INJECT1_1 = "NO";
    LUT4 i7_4_lut (.A(\spi_cmd_r[7] ), .B(\spi_cmd_r[10] ), .C(spi_data_valid_r), 
         .D(\spi_cmd_r[12] ), .Z(n18)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i7_4_lut.init = 16'h0010;
    CCU2D equal_10_13 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24935), 
          .S0(pwm_N_898));
    defparam equal_10_13.INIT0 = 16'hFFFF;
    defparam equal_10_13.INIT1 = 16'h0000;
    defparam equal_10_13.INJECT1_0 = "NO";
    defparam equal_10_13.INJECT1_1 = "NO";
    CCU2D equal_10_9 (.A0(pwm_N_899[11]), .B0(pwm_freq_cntr[11]), .C0(pwm_N_899[10]), 
          .D0(pwm_freq_cntr[10]), .A1(pwm_N_899[9]), .B1(pwm_freq_cntr[9]), 
          .C1(pwm_N_899[8]), .D1(pwm_freq_cntr[8]), .CIN(n24932), .COUT(n24933));
    defparam equal_10_9.INIT0 = 16'h9009;
    defparam equal_10_9.INIT1 = 16'h9009;
    defparam equal_10_9.INJECT1_0 = "YES";
    defparam equal_10_9.INJECT1_1 = "YES";
    CCU2D equal_10_13_20020 (.A0(pwm_N_899[3]), .B0(pwm_freq_cntr[3]), .C0(pwm_N_899[2]), 
          .D0(pwm_freq_cntr[2]), .A1(pwm_N_899[1]), .B1(pwm_freq_cntr[1]), 
          .C1(pwm_N_899[0]), .D1(pwm_freq_cntr[0]), .CIN(n24934), .COUT(n24935));
    defparam equal_10_13_20020.INIT0 = 16'h9009;
    defparam equal_10_13_20020.INIT1 = 16'h9009;
    defparam equal_10_13_20020.INJECT1_0 = "YES";
    defparam equal_10_13_20020.INJECT1_1 = "YES";
    CCU2D pwm_freq_cntr_2503_add_4_13 (.A0(pwm_freq_cntr[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25205), .S0(n53[11]));   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503_add_4_13.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_2503_add_4_13.INIT1 = 16'h0000;
    defparam pwm_freq_cntr_2503_add_4_13.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_2503_add_4_13.INJECT1_1 = "NO";
    CCU2D add_395_3 (.A0(status_cntr[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(status_cntr[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24968), .COUT(n24969), .S0(n827[1]), .S1(n827[2]));   // c:/s_links/sources/status_led.v(59[19:34])
    defparam add_395_3.INIT0 = 16'h5aaa;
    defparam add_395_3.INIT1 = 16'h5aaa;
    defparam add_395_3.INJECT1_0 = "NO";
    defparam add_395_3.INJECT1_1 = "NO";
    CCU2D add_395_11 (.A0(status_cntr[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(status_cntr[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24972), .COUT(n24973), .S0(n827[9]), .S1(n827[10]));   // c:/s_links/sources/status_led.v(59[19:34])
    defparam add_395_11.INIT0 = 16'h5aaa;
    defparam add_395_11.INIT1 = 16'h5aaa;
    defparam add_395_11.INJECT1_0 = "NO";
    defparam add_395_11.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_2503_add_4_11 (.A0(pwm_freq_cntr[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[10]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n25204), .COUT(n25205), .S0(n53[9]), 
          .S1(n53[10]));   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503_add_4_11.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_2503_add_4_11.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_2503_add_4_11.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_2503_add_4_11.INJECT1_1 = "NO";
    LUT4 i22444_2_lut (.A(\spi_cmd_r[6] ), .B(\spi_cmd_r[15] ), .Z(n27614)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22444_2_lut.init = 16'heeee;
    CCU2D pwm_freq_cntr_2503_add_4_9 (.A0(pwm_freq_cntr[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[8]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n25203), .COUT(n25204), .S0(n53[7]), 
          .S1(n53[8]));   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503_add_4_9.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_2503_add_4_9.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_2503_add_4_9.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_2503_add_4_9.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_2503_add_4_7 (.A0(pwm_freq_cntr[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n25202), .COUT(n25203), .S0(n53[5]), 
          .S1(n53[6]));   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503_add_4_7.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_2503_add_4_7.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_2503_add_4_7.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_2503_add_4_7.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_2503_add_4_5 (.A0(pwm_freq_cntr[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n25201), .COUT(n25202), .S0(n53[3]), 
          .S1(n53[4]));   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503_add_4_5.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_2503_add_4_5.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_2503_add_4_5.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_2503_add_4_5.INJECT1_1 = "NO";
    CCU2D pwm_freq_cntr_2503_add_4_3 (.A0(pwm_freq_cntr[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(pwm_freq_cntr[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n25200), .COUT(n25201), .S0(n53[1]), 
          .S1(n53[2]));   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503_add_4_3.INIT0 = 16'hfaaa;
    defparam pwm_freq_cntr_2503_add_4_3.INIT1 = 16'hfaaa;
    defparam pwm_freq_cntr_2503_add_4_3.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_2503_add_4_3.INJECT1_1 = "NO";
    LUT4 i1_3_lut (.A(pwm_N_898), .B(resetn_c), .C(n14283), .Z(clk_enable_517)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i1_3_lut.init = 16'hc8c8;
    CCU2D pwm_freq_cntr_2503_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_freq_cntr[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n25200), .S1(n53[0]));   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503_add_4_1.INIT0 = 16'hF000;
    defparam pwm_freq_cntr_2503_add_4_1.INIT1 = 16'h0555;
    defparam pwm_freq_cntr_2503_add_4_1.INJECT1_0 = "NO";
    defparam pwm_freq_cntr_2503_add_4_1.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_13 (.A0(pwm_duty[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25050), .S0(pwm_N_899[11]), .S1(pwm_N_899[12]));   // c:/s_links/sources/status_led.v(66[29:41])
    defparam sub_14_add_2_13.INIT0 = 16'h5555;
    defparam sub_14_add_2_13.INIT1 = 16'hffff;
    defparam sub_14_add_2_13.INJECT1_0 = "NO";
    defparam sub_14_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_11 (.A0(pwm_duty[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25049), .COUT(n25050), .S0(pwm_N_899[9]), 
          .S1(pwm_N_899[10]));   // c:/s_links/sources/status_led.v(66[29:41])
    defparam sub_14_add_2_11.INIT0 = 16'h5555;
    defparam sub_14_add_2_11.INIT1 = 16'h5555;
    defparam sub_14_add_2_11.INJECT1_0 = "NO";
    defparam sub_14_add_2_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(n14283), .B(n17), .C(n22), .D(n18_adj_7606), .Z(pwm_N_896)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut.init = 16'haaa8;
    CCU2D sub_14_add_2_9 (.A0(pwm_duty[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25048), .COUT(n25049), .S0(pwm_N_899[7]), 
          .S1(pwm_N_899[8]));   // c:/s_links/sources/status_led.v(66[29:41])
    defparam sub_14_add_2_9.INIT0 = 16'h5555;
    defparam sub_14_add_2_9.INIT1 = 16'h5555;
    defparam sub_14_add_2_9.INJECT1_0 = "NO";
    defparam sub_14_add_2_9.INJECT1_1 = "NO";
    LUT4 i5_2_lut (.A(pwm_duty[4]), .B(pwm_duty[7]), .Z(n17)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/status_led.v(61[8:23])
    defparam i5_2_lut.init = 16'heeee;
    CCU2D sub_14_add_2_7 (.A0(pwm_duty[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25047), .COUT(n25048), .S0(pwm_N_899[5]), 
          .S1(pwm_N_899[6]));   // c:/s_links/sources/status_led.v(66[29:41])
    defparam sub_14_add_2_7.INIT0 = 16'h5555;
    defparam sub_14_add_2_7.INIT1 = 16'h5555;
    defparam sub_14_add_2_7.INJECT1_0 = "NO";
    defparam sub_14_add_2_7.INJECT1_1 = "NO";
    LUT4 i10_4_lut_adj_956 (.A(pwm_duty[10]), .B(n20), .C(n14_adj_7607), 
         .D(pwm_duty[0]), .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/status_led.v(61[8:23])
    defparam i10_4_lut_adj_956.init = 16'hfffe;
    CCU2D sub_14_add_2_5 (.A0(pwm_duty[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25046), .COUT(n25047), .S0(pwm_N_899[3]), 
          .S1(pwm_N_899[4]));   // c:/s_links/sources/status_led.v(66[29:41])
    defparam sub_14_add_2_5.INIT0 = 16'h5555;
    defparam sub_14_add_2_5.INIT1 = 16'h5555;
    defparam sub_14_add_2_5.INJECT1_0 = "NO";
    defparam sub_14_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_3 (.A0(pwm_duty[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pwm_duty[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25045), .COUT(n25046), .S0(pwm_N_899[1]), 
          .S1(pwm_N_899[2]));   // c:/s_links/sources/status_led.v(66[29:41])
    defparam sub_14_add_2_3.INIT0 = 16'h5555;
    defparam sub_14_add_2_3.INIT1 = 16'h5555;
    defparam sub_14_add_2_3.INJECT1_0 = "NO";
    defparam sub_14_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_14_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_duty[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n25045), .S1(pwm_N_899[0]));   // c:/s_links/sources/status_led.v(66[29:41])
    defparam sub_14_add_2_1.INIT0 = 16'hF000;
    defparam sub_14_add_2_1.INIT1 = 16'h5555;
    defparam sub_14_add_2_1.INJECT1_0 = "NO";
    defparam sub_14_add_2_1.INJECT1_1 = "NO";
    LUT4 i6_2_lut (.A(pwm_duty[1]), .B(pwm_duty[2]), .Z(n18_adj_7606)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/status_led.v(61[8:23])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i8_4_lut_adj_957 (.A(pwm_duty[9]), .B(pwm_duty[6]), .C(pwm_duty[3]), 
         .D(pwm_duty[11]), .Z(n20)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/status_led.v(61[8:23])
    defparam i8_4_lut_adj_957.init = 16'hfffe;
    LUT4 i2_2_lut (.A(pwm_duty[5]), .B(pwm_duty[8]), .Z(n14_adj_7607)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/status_led.v(61[8:23])
    defparam i2_2_lut.init = 16'heeee;
    CCU2D equal_10_11 (.A0(pwm_N_899[7]), .B0(pwm_freq_cntr[7]), .C0(pwm_N_899[6]), 
          .D0(pwm_freq_cntr[6]), .A1(pwm_N_899[5]), .B1(pwm_freq_cntr[5]), 
          .C1(pwm_N_899[4]), .D1(pwm_freq_cntr[4]), .CIN(n24933), .COUT(n24934));
    defparam equal_10_11.INIT0 = 16'h9009;
    defparam equal_10_11.INIT1 = 16'h9009;
    defparam equal_10_11.INJECT1_0 = "YES";
    defparam equal_10_11.INJECT1_1 = "YES";
    CCU2D add_395_5 (.A0(status_cntr[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(status_cntr[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24969), .COUT(n24970), .S0(n827[3]), .S1(n827[4]));   // c:/s_links/sources/status_led.v(59[19:34])
    defparam add_395_5.INIT0 = 16'h5aaa;
    defparam add_395_5.INIT1 = 16'h5aaa;
    defparam add_395_5.INJECT1_0 = "NO";
    defparam add_395_5.INJECT1_1 = "NO";
    CCU2D add_395_13 (.A0(status_cntr[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(status_cntr[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n24973), .S0(n827[11]), .S1(n827[12]));   // c:/s_links/sources/status_led.v(59[19:34])
    defparam add_395_13.INIT0 = 16'h5aaa;
    defparam add_395_13.INIT1 = 16'h5aaa;
    defparam add_395_13.INJECT1_0 = "NO";
    defparam add_395_13.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_491 (.A(status_cntr[10]), .B(status_cntr[9]), .C(status_cntr[8]), 
         .Z(n29219)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut_rep_491.init = 16'h8080;
    LUT4 i1_2_lut_4_lut (.A(status_cntr[10]), .B(status_cntr[9]), .C(status_cntr[8]), 
         .D(status_cntr[7]), .Z(n26939)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_adj_958 (.A(n14283), .B(n827[6]), .Z(n141[6])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_958.init = 16'h8888;
    FD1P3IX pwm_duty__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_303), .CD(n29239), 
            .CK(clk), .Q(pwm_duty[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i11.GSR = "DISABLED";
    FD1P3IX pwm_duty__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_303), .CD(n29239), 
            .CK(clk), .Q(pwm_duty[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i10.GSR = "DISABLED";
    FD1P3IX pwm_duty__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_303), .CD(n29239), 
            .CK(clk), .Q(pwm_duty[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i9.GSR = "DISABLED";
    FD1P3IX pwm_duty__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_303), .CD(n29239), 
            .CK(clk), .Q(pwm_duty[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i8.GSR = "DISABLED";
    FD1P3IX pwm_duty__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_303), .CD(n29239), 
            .CK(clk), .Q(pwm_duty[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i7.GSR = "DISABLED";
    FD1P3IX pwm_duty__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_303), .CD(n29239), 
            .CK(clk), .Q(pwm_duty[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i6.GSR = "DISABLED";
    FD1P3IX pwm_duty__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_303), .CD(n29239), 
            .CK(clk), .Q(pwm_duty[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i5.GSR = "DISABLED";
    FD1P3IX pwm_duty__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_303), .CD(n29239), 
            .CK(clk), .Q(pwm_duty[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i4.GSR = "DISABLED";
    FD1P3IX pwm_duty__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_303), .CD(n29239), 
            .CK(clk), .Q(pwm_duty[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i3.GSR = "DISABLED";
    FD1P3IX pwm_duty__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_303), .CD(n29239), 
            .CK(clk), .Q(pwm_duty[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i2.GSR = "DISABLED";
    FD1P3IX pwm_duty__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_303), .CD(n29239), 
            .CK(clk), .Q(pwm_duty[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_duty__i1.GSR = "DISABLED";
    FD1P3IX status_cntr_i0_i0 (.D(n827[0]), .SP(clk_enable_308), .CD(n14229), 
            .CK(clk), .Q(status_cntr[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam status_cntr_i0_i0.GSR = "DISABLED";
    LUT4 i1_2_lut_adj_959 (.A(n14283), .B(n827[7]), .Z(n141[7])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_959.init = 16'h8888;
    LUT4 i14662_4_lut_rep_385 (.A(n29755), .B(resetn_c), .C(n14283), .D(n6), 
         .Z(clk_enable_308)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i14662_4_lut_rep_385.init = 16'hccc8;
    LUT4 i1_2_lut_adj_960 (.A(n14283), .B(n827[8]), .Z(n141[8])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_960.init = 16'h8888;
    LUT4 i5_3_lut_adj_961 (.A(\spi_addr[3] ), .B(n10), .C(n27465), .Z(n13490)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i5_3_lut_adj_961.init = 16'hfdfd;
    LUT4 i1_2_lut_adj_962 (.A(n14283), .B(n827[9]), .Z(n141[9])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_962.init = 16'h8888;
    LUT4 i4_4_lut (.A(\spi_cmd[1] ), .B(\spi_addr[0] ), .C(n13489), .D(n26928), 
         .Z(n10)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i4_4_lut.init = 16'hfffb;
    LUT4 i1_2_lut_adj_963 (.A(n14283), .B(n827[10]), .Z(n141[10])) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_963.init = 16'h8888;
    FD1P3AX pwm_341 (.D(pwm_N_896), .SP(clk_enable_517), .CK(clk), .Q(pwm)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=228, LSE_RLINE=245 */ ;   // c:/s_links/sources/status_led.v(40[8] 92[4])
    defparam pwm_341.GSR = "DISABLED";
    LUT4 i1_2_lut_adj_964 (.A(n14160), .B(status_cntr[12]), .Z(pwm_out_N_893)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_964.init = 16'heeee;
    LUT4 i9206_4_lut (.A(n26939), .B(status_cntr[11]), .C(status_cntr[6]), 
         .D(n12), .Z(n14160)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i9206_4_lut.init = 16'heccc;
    LUT4 i3348_2_lut (.A(status_cntr[4]), .B(status_cntr[5]), .Z(n12)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3348_2_lut.init = 16'heeee;
    LUT4 i22589_3_lut (.A(n19475), .B(resetn_c), .C(status_cntr[12]), 
         .Z(clk_enable_205)) /* synthesis lut_function=(!(A (B (C)))) */ ;
    defparam i22589_3_lut.init = 16'h7f7f;
    LUT4 i1_3_lut_adj_965 (.A(resetn_c), .B(n14161), .C(status_cntr[12]), 
         .Z(n27015)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i1_3_lut_adj_965.init = 16'h0808;
    LUT4 i9207_4_lut (.A(pwm), .B(n26939), .C(n14160), .D(n4), .Z(n14161)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B ((D)+!C)+!B !(C)))) */ ;   // c:/s_links/sources/status_led.v(87[8] 90[6])
    defparam i9207_4_lut.init = 16'h3afa;
    LUT4 i1_3_lut_adj_966 (.A(status_cntr[5]), .B(status_cntr[11]), .C(status_cntr[6]), 
         .Z(n4)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i1_3_lut_adj_966.init = 16'hc8c8;
    LUT4 i14535_4_lut (.A(n25288), .B(status_cntr[11]), .C(n29219), .D(status_cntr[7]), 
         .Z(n19475)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i14535_4_lut.init = 16'hfcec;
    LUT4 i2_3_lut (.A(status_cntr[6]), .B(status_cntr[4]), .C(status_cntr[5]), 
         .Z(n25288)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    CCU2D equal_10_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(pwm_N_899[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24932));   // c:/s_links/sources/status_led.v(66[12:41])
    defparam equal_10_0.INIT0 = 16'hF000;
    defparam equal_10_0.INIT1 = 16'h5555;
    defparam equal_10_0.INJECT1_0 = "NO";
    defparam equal_10_0.INJECT1_1 = "YES";
    FD1P3IX pwm_freq_cntr_2503__i11 (.D(n53[11]), .SP(resetn_c), .CD(n14284), 
            .CK(clk), .Q(pwm_freq_cntr[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503__i11.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_2503__i10 (.D(n53[10]), .SP(resetn_c), .CD(n14284), 
            .CK(clk), .Q(pwm_freq_cntr[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503__i10.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_2503__i9 (.D(n53[9]), .SP(resetn_c), .CD(n14284), 
            .CK(clk), .Q(pwm_freq_cntr[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503__i9.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_2503__i8 (.D(n53[8]), .SP(resetn_c), .CD(n14284), 
            .CK(clk), .Q(pwm_freq_cntr[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503__i8.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_2503__i7 (.D(n53[7]), .SP(resetn_c), .CD(n14284), 
            .CK(clk), .Q(pwm_freq_cntr[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503__i7.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_2503__i6 (.D(n53[6]), .SP(resetn_c), .CD(n14284), 
            .CK(clk), .Q(pwm_freq_cntr[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503__i6.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_2503__i5 (.D(n53[5]), .SP(resetn_c), .CD(n14284), 
            .CK(clk), .Q(pwm_freq_cntr[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503__i5.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_2503__i4 (.D(n53[4]), .SP(resetn_c), .CD(n14284), 
            .CK(clk), .Q(pwm_freq_cntr[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503__i4.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_2503__i3 (.D(n53[3]), .SP(resetn_c), .CD(n14284), 
            .CK(clk), .Q(pwm_freq_cntr[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503__i3.GSR = "DISABLED";
    FD1P3IX pwm_freq_cntr_2503__i2 (.D(n53[2]), .SP(resetn_c), .CD(n14284), 
            .CK(clk), .Q(pwm_freq_cntr[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/status_led.v(71[22:42])
    defparam pwm_freq_cntr_2503__i2.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \intrpt_ctrl(DEV_ID=4) 
//

module \intrpt_ctrl(DEV_ID=4)  (\spi_data_out_r_39__N_2856[0] , clk, \pin_intrpt[12] , 
            n29239, clear_intrpt, clear_intrpt_N_2923, intrpt_out_c_4, 
            intrpt_out_N_2919, n29757, \spi_data_out_r_39__N_2856[2] , 
            \pin_intrpt[14] , \spi_data_out_r_39__N_2856[1] , \pin_intrpt[13] ) /* synthesis syn_module_defined=1 */ ;
    output \spi_data_out_r_39__N_2856[0] ;
    input clk;
    input \pin_intrpt[12] ;
    input n29239;
    output clear_intrpt;
    input clear_intrpt_N_2923;
    output intrpt_out_c_4;
    input intrpt_out_N_2919;
    input n29757;
    output \spi_data_out_r_39__N_2856[2] ;
    input \pin_intrpt[14] ;
    output \spi_data_out_r_39__N_2856[1] ;
    input \pin_intrpt[13] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire \pin_intrpt[14]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[14] */ ;   // c:/s_links/sources/mcm_top.v(102[46:56])
    wire [2:0]intrpt_in_reg;   // c:/s_links/sources/intrpt_ctrl.v(38[35:48])
    wire [2:0]intrpt_in_dly;   // c:/s_links/sources/intrpt_ctrl.v(39[36:49])
    
    wire assert_intrpt, intrpt_all_edges, n4;
    
    FD1S3AX spi_data_out_r_i1 (.D(\pin_intrpt[12] ), .CK(clk), .Q(\spi_data_out_r_39__N_2856[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i0 (.D(\pin_intrpt[12] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i0.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i0 (.D(intrpt_in_reg[0]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i0.GSR = "DISABLED";
    FD1S3IX clear_intrpt_317 (.D(clear_intrpt_N_2923), .CK(clk), .CD(n29239), 
            .Q(clear_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam clear_intrpt_317.GSR = "DISABLED";
    FD1S3IX assert_intrpt_316 (.D(intrpt_all_edges), .CK(clk), .CD(n29239), 
            .Q(assert_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(63[8] 73[4])
    defparam assert_intrpt_316.GSR = "DISABLED";
    FD1P3IX intrpt_out_359 (.D(n29757), .SP(assert_intrpt), .CD(intrpt_out_N_2919), 
            .CK(clk), .Q(intrpt_out_c_4)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(92[8] 99[4])
    defparam intrpt_out_359.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\pin_intrpt[14] ), .CK(clk), .Q(\spi_data_out_r_39__N_2856[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\pin_intrpt[13] ), .CK(clk), .Q(\spi_data_out_r_39__N_2856[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i1 (.D(\pin_intrpt[13] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i2 (.D(\pin_intrpt[14] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i1 (.D(intrpt_in_reg[1]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i2 (.D(intrpt_in_reg[2]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i2.GSR = "DISABLED";
    LUT4 i2_3_lut (.A(intrpt_in_dly[0]), .B(n4), .C(intrpt_in_reg[0]), 
         .Z(intrpt_all_edges)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i2_3_lut.init = 16'hdede;
    LUT4 i1_4_lut (.A(intrpt_in_dly[1]), .B(intrpt_in_dly[2]), .C(intrpt_in_reg[1]), 
         .D(intrpt_in_reg[2]), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i1_4_lut.init = 16'h7bde;
    
endmodule
//
// Verilog Description of module \intrpt_ctrl(DEV_ID=3) 
//

module \intrpt_ctrl(DEV_ID=3)  (clk, n29239, \spi_data_out_r_39__N_2785[0] , 
            \pin_intrpt[9] , clear_intrpt, clear_intrpt_N_2852, intrpt_out_c_3, 
            intrpt_out_N_2848, n29757, \spi_data_out_r_39__N_2785[2] , 
            \pin_intrpt[11] , \spi_data_out_r_39__N_2785[1] , \pin_intrpt[10] ) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input n29239;
    output \spi_data_out_r_39__N_2785[0] ;
    input \pin_intrpt[9] ;
    output clear_intrpt;
    input clear_intrpt_N_2852;
    output intrpt_out_c_3;
    input intrpt_out_N_2848;
    input n29757;
    output \spi_data_out_r_39__N_2785[2] ;
    input \pin_intrpt[11] ;
    output \spi_data_out_r_39__N_2785[1] ;
    input \pin_intrpt[10] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire \pin_intrpt[11]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[11] */ ;   // c:/s_links/sources/mcm_top.v(102[46:56])
    wire [2:0]intrpt_in_dly;   // c:/s_links/sources/intrpt_ctrl.v(39[36:49])
    wire [2:0]intrpt_in_reg;   // c:/s_links/sources/intrpt_ctrl.v(38[35:48])
    
    wire assert_intrpt, intrpt_all_edges, n4;
    
    FD1S3IX intrpt_in_dly__i0 (.D(intrpt_in_reg[0]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\pin_intrpt[9] ), .CK(clk), .Q(\spi_data_out_r_39__N_2785[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i0 (.D(\pin_intrpt[9] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i0.GSR = "DISABLED";
    FD1S3IX clear_intrpt_317 (.D(clear_intrpt_N_2852), .CK(clk), .CD(n29239), 
            .Q(clear_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam clear_intrpt_317.GSR = "DISABLED";
    FD1S3IX assert_intrpt_316 (.D(intrpt_all_edges), .CK(clk), .CD(n29239), 
            .Q(assert_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(63[8] 73[4])
    defparam assert_intrpt_316.GSR = "DISABLED";
    FD1P3IX intrpt_out_359 (.D(n29757), .SP(assert_intrpt), .CD(intrpt_out_N_2848), 
            .CK(clk), .Q(intrpt_out_c_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(92[8] 99[4])
    defparam intrpt_out_359.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\pin_intrpt[11] ), .CK(clk), .Q(\spi_data_out_r_39__N_2785[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\pin_intrpt[10] ), .CK(clk), .Q(\spi_data_out_r_39__N_2785[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i2 (.D(intrpt_in_reg[2]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i1 (.D(intrpt_in_reg[1]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i1 (.D(\pin_intrpt[10] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i2 (.D(\pin_intrpt[11] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i2.GSR = "DISABLED";
    LUT4 i2_3_lut (.A(intrpt_in_dly[0]), .B(n4), .C(intrpt_in_reg[0]), 
         .Z(intrpt_all_edges)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i2_3_lut.init = 16'hdede;
    LUT4 i1_4_lut (.A(intrpt_in_dly[1]), .B(intrpt_in_dly[2]), .C(intrpt_in_reg[1]), 
         .D(intrpt_in_reg[2]), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i1_4_lut.init = 16'h7bde;
    
endmodule
//
// Verilog Description of module \intrpt_ctrl(DEV_ID=2) 
//

module \intrpt_ctrl(DEV_ID=2)  (clk, n29239, \spi_data_out_r_39__N_2714[0] , 
            \pin_intrpt[6] , intrpt_out_c_2, intrpt_out_N_2777, n29757, 
            clear_intrpt, clear_intrpt_N_2781, \spi_data_out_r_39__N_2714[2] , 
            \mode[2]_derived_32 , \spi_data_out_r_39__N_2714[1] , \pin_intrpt[7] ) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input n29239;
    output \spi_data_out_r_39__N_2714[0] ;
    input \pin_intrpt[6] ;
    output intrpt_out_c_2;
    input intrpt_out_N_2777;
    input n29757;
    output clear_intrpt;
    input clear_intrpt_N_2781;
    output \spi_data_out_r_39__N_2714[2] ;
    input \mode[2]_derived_32 ;
    output \spi_data_out_r_39__N_2714[1] ;
    input \pin_intrpt[7] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire \mode[2]_derived_32  /* synthesis is_clock=1, SET_AS_NETWORK=\stepper_ins[2].u_stepper/mode[2]_derived_32 */ ;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    wire [2:0]intrpt_in_dly;   // c:/s_links/sources/intrpt_ctrl.v(39[36:49])
    wire [2:0]intrpt_in_reg;   // c:/s_links/sources/intrpt_ctrl.v(38[35:48])
    
    wire assert_intrpt, intrpt_all_edges, n4;
    
    FD1S3IX intrpt_in_dly__i0 (.D(intrpt_in_reg[0]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\pin_intrpt[6] ), .CK(clk), .Q(\spi_data_out_r_39__N_2714[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i0 (.D(\pin_intrpt[6] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i0.GSR = "DISABLED";
    FD1P3IX intrpt_out_359 (.D(n29757), .SP(assert_intrpt), .CD(intrpt_out_N_2777), 
            .CK(clk), .Q(intrpt_out_c_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(92[8] 99[4])
    defparam intrpt_out_359.GSR = "DISABLED";
    FD1S3IX clear_intrpt_317 (.D(clear_intrpt_N_2781), .CK(clk), .CD(n29239), 
            .Q(clear_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam clear_intrpt_317.GSR = "DISABLED";
    FD1S3IX assert_intrpt_316 (.D(intrpt_all_edges), .CK(clk), .CD(n29239), 
            .Q(assert_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(63[8] 73[4])
    defparam assert_intrpt_316.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\mode[2]_derived_32 ), .CK(clk), .Q(\spi_data_out_r_39__N_2714[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\pin_intrpt[7] ), .CK(clk), .Q(\spi_data_out_r_39__N_2714[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i2 (.D(intrpt_in_reg[2]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i1 (.D(intrpt_in_reg[1]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i1 (.D(\pin_intrpt[7] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i2 (.D(\mode[2]_derived_32 ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i2.GSR = "DISABLED";
    LUT4 i2_3_lut (.A(intrpt_in_dly[0]), .B(n4), .C(intrpt_in_reg[0]), 
         .Z(intrpt_all_edges)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i2_3_lut.init = 16'hdede;
    LUT4 i1_4_lut (.A(intrpt_in_dly[1]), .B(intrpt_in_dly[2]), .C(intrpt_in_reg[1]), 
         .D(intrpt_in_reg[2]), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i1_4_lut.init = 16'h7bde;
    
endmodule
//
// Verilog Description of module cs_decoder
//

module cs_decoder (cs_decoded, CS_READY_c, FLASH_CS_c, MAX3421_CS_c, 
            cs_c_0, cs_c_1, cs_c_2, cs_c_4, cs_c_3) /* synthesis syn_module_defined=1 */ ;
    output [13:0]cs_decoded;
    input CS_READY_c;
    output FLASH_CS_c;
    output MAX3421_CS_c;
    input cs_c_0;
    input cs_c_1;
    input cs_c_2;
    input cs_c_4;
    input cs_c_3;
    
    wire CS_READY_c /* synthesis is_clock=1, SET_AS_NETWORK=CS_READY_c */ ;   // c:/s_links/sources/mcm_top.v(23[24:32])
    
    wire CS_READY_c_enable_1;
    wire [13:0]cs_decoded_13__N_752;
    
    wire CS_READY_c_enable_2, FLASH_CS_N_768, CS_READY_c_enable_3, CS_READY_c_enable_4, 
        CS_READY_c_enable_5, CS_READY_c_enable_6, n28852, n29236, n33, 
        n29330, n29331, n29133, n10262, n29258, n29292, n13889, 
        n29197, n29274, n29163, CS_READY_c_enable_14, n29188, n29131, 
        n29272, n29273, n29159, n71, n27352, CS_READY_c_enable_7, 
        CS_READY_c_enable_8, CS_READY_c_enable_9, CS_READY_c_enable_10, 
        CS_READY_c_enable_11, CS_READY_c_enable_12, CS_READY_c_enable_13, 
        CS_READY_c_enable_15, CS_READY_c_enable_16, n27728, n27736, 
        n27513;
    
    FD1P3AY cs_decoded_i0 (.D(cs_decoded_13__N_752[0]), .SP(CS_READY_c_enable_1), 
            .CK(CS_READY_c), .Q(cs_decoded[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i0.GSR = "ENABLED";
    FD1P3AY FLASH_CS_14 (.D(FLASH_CS_N_768), .SP(CS_READY_c_enable_2), .CK(CS_READY_c), 
            .Q(FLASH_CS_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam FLASH_CS_14.GSR = "ENABLED";
    FD1P3AY MAX3421_CS_15 (.D(FLASH_CS_N_768), .SP(CS_READY_c_enable_3), 
            .CK(CS_READY_c), .Q(MAX3421_CS_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam MAX3421_CS_15.GSR = "ENABLED";
    FD1P3AY cs_decoded_i1 (.D(cs_decoded_13__N_752[2]), .SP(CS_READY_c_enable_4), 
            .CK(CS_READY_c), .Q(cs_decoded[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i1.GSR = "ENABLED";
    FD1P3AY cs_decoded_i2 (.D(cs_decoded_13__N_752[2]), .SP(CS_READY_c_enable_5), 
            .CK(CS_READY_c), .Q(cs_decoded[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i2.GSR = "ENABLED";
    FD1P3AY cs_decoded_i3 (.D(cs_decoded_13__N_752[3]), .SP(CS_READY_c_enable_6), 
            .CK(CS_READY_c), .Q(cs_decoded[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i3.GSR = "ENABLED";
    LUT4 n28852_bdd_2_lut (.A(n28852), .B(cs_c_0), .Z(CS_READY_c_enable_3)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n28852_bdd_2_lut.init = 16'h2222;
    LUT4 i22567_2_lut_rep_508 (.A(cs_c_1), .B(cs_c_0), .Z(n29236)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i22567_2_lut_rep_508.init = 16'h6666;
    LUT4 i1_2_lut_3_lut (.A(cs_c_1), .B(cs_c_0), .C(cs_c_2), .Z(n33)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+(C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h0909;
    PFUMX i23162 (.BLUT(n29330), .ALUT(n29331), .C0(cs_c_4), .Z(CS_READY_c_enable_2));
    LUT4 i2_4_lut (.A(cs_c_3), .B(n29133), .C(cs_c_4), .D(n10262), .Z(CS_READY_c_enable_1)) /* synthesis lut_function=(A (B)+!A (B (C+!(D)))) */ ;
    defparam i2_4_lut.init = 16'hc8cc;
    LUT4 i5469_2_lut (.A(cs_c_1), .B(cs_c_2), .Z(n10262)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/cs_decoder.v(32[5] 74[10])
    defparam i5469_2_lut.init = 16'heeee;
    LUT4 i111_2_lut_rep_530 (.A(cs_c_0), .B(cs_c_2), .Z(n29258)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i111_2_lut_rep_530.init = 16'heeee;
    LUT4 i1_3_lut_4_lut (.A(cs_c_0), .B(cs_c_2), .C(n29292), .D(cs_c_1), 
         .Z(n13889)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i2_3_lut_4_lut_4_lut (.A(n29197), .B(n29274), .C(n13889), .D(n29163), 
         .Z(CS_READY_c_enable_14)) /* synthesis lut_function=(!(A (D)+!A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i2_3_lut_4_lut_4_lut.init = 16'h00ea;
    LUT4 i1_2_lut_rep_403_3_lut (.A(n29188), .B(cs_c_4), .C(n13889), .Z(n29131)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam i1_2_lut_rep_403_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_544 (.A(cs_c_2), .B(cs_c_3), .Z(n29272)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_2_lut_rep_544.init = 16'h8888;
    LUT4 i1_3_lut_rep_460_4_lut (.A(cs_c_2), .B(cs_c_3), .C(cs_c_1), .D(cs_c_0), 
         .Z(n29188)) /* synthesis lut_function=(!(((C (D)+!C !(D))+!B)+!A)) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_3_lut_rep_460_4_lut.init = 16'h0880;
    LUT4 i1_2_lut_rep_545 (.A(cs_c_0), .B(cs_c_2), .Z(n29273)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_2_lut_rep_545.init = 16'h8888;
    LUT4 i1_2_lut_rep_431_3_lut_4_lut (.A(cs_c_0), .B(cs_c_2), .C(n29274), 
         .D(cs_c_1), .Z(n29159)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_2_lut_rep_431_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i79_3_lut_4_lut_3_lut (.A(cs_c_0), .B(cs_c_2), .C(cs_c_1), .Z(n71)) /* synthesis lut_function=(A (B (C))+!A !(B+(C))) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i79_3_lut_4_lut_3_lut.init = 16'h8181;
    LUT4 i1_2_lut_rep_469_3_lut (.A(cs_c_0), .B(cs_c_2), .C(cs_c_1), .Z(n29197)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_2_lut_rep_469_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_546 (.A(cs_c_4), .B(cs_c_3), .Z(n29274)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_2_lut_rep_546.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_adj_946 (.A(cs_c_4), .B(cs_c_3), .C(cs_c_0), .Z(cs_decoded_13__N_752[13])) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_2_lut_3_lut_adj_946.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_947 (.A(cs_c_4), .B(cs_c_3), .C(cs_c_1), .Z(cs_decoded_13__N_752[12])) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_2_lut_3_lut_adj_947.init = 16'hfbfb;
    LUT4 i1_2_lut_rep_405_3_lut_4_lut_4_lut (.A(cs_c_4), .B(cs_c_3), .C(n29197), 
         .D(n29188), .Z(n29133)) /* synthesis lut_function=(!(A (D)+!A !((C)+!B))) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_2_lut_rep_405_3_lut_4_lut_4_lut.init = 16'h51fb;
    LUT4 i9125_2_lut_rep_435_4_lut (.A(cs_c_0), .B(n29272), .C(cs_c_1), 
         .D(cs_c_4), .Z(n29163)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C (D))))) */ ;   // c:/s_links/sources/cs_decoder.v(32[5] 74[10])
    defparam i9125_2_lut_rep_435_4_lut.init = 16'h4800;
    LUT4 i1_2_lut_3_lut_adj_948 (.A(cs_c_4), .B(cs_c_3), .C(cs_c_2), .Z(cs_decoded_13__N_752[9])) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_2_lut_3_lut_adj_948.init = 16'hfbfb;
    LUT4 i1_3_lut_4_lut_adj_949 (.A(cs_c_1), .B(n29273), .C(cs_c_3), .D(cs_c_4), 
         .Z(n27352)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_3_lut_4_lut_adj_949.init = 16'hff80;
    LUT4 i1_2_lut_rep_564 (.A(cs_c_3), .B(cs_c_4), .Z(n29292)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_2_lut_rep_564.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_950 (.A(cs_c_3), .B(cs_c_4), .C(cs_c_0), .Z(cs_decoded_13__N_752[0])) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_2_lut_3_lut_adj_950.init = 16'hefef;
    LUT4 i1_2_lut_3_lut_adj_951 (.A(cs_c_3), .B(cs_c_4), .C(cs_c_2), .Z(cs_decoded_13__N_752[6])) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_2_lut_3_lut_adj_951.init = 16'hefef;
    FD1P3AY cs_decoded_i13 (.D(cs_decoded_13__N_752[13]), .SP(CS_READY_c_enable_7), 
            .CK(CS_READY_c), .Q(cs_decoded[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i13.GSR = "ENABLED";
    FD1P3AY cs_decoded_i12 (.D(cs_decoded_13__N_752[12]), .SP(CS_READY_c_enable_8), 
            .CK(CS_READY_c), .Q(cs_decoded[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i12.GSR = "ENABLED";
    FD1P3AY cs_decoded_i11 (.D(cs_decoded_13__N_752[12]), .SP(CS_READY_c_enable_9), 
            .CK(CS_READY_c), .Q(cs_decoded[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i11.GSR = "ENABLED";
    FD1P3AY cs_decoded_i10 (.D(cs_decoded_13__N_752[9]), .SP(CS_READY_c_enable_10), 
            .CK(CS_READY_c), .Q(cs_decoded[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i10.GSR = "ENABLED";
    FD1P3AY cs_decoded_i9 (.D(cs_decoded_13__N_752[9]), .SP(CS_READY_c_enable_11), 
            .CK(CS_READY_c), .Q(cs_decoded[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i9.GSR = "ENABLED";
    FD1P3AY cs_decoded_i8 (.D(cs_decoded_13__N_752[9]), .SP(CS_READY_c_enable_12), 
            .CK(CS_READY_c), .Q(cs_decoded[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i8.GSR = "ENABLED";
    FD1P3AY cs_decoded_i7 (.D(cs_decoded_13__N_752[9]), .SP(CS_READY_c_enable_13), 
            .CK(CS_READY_c), .Q(cs_decoded[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i7.GSR = "ENABLED";
    FD1P3AY cs_decoded_i6 (.D(cs_decoded_13__N_752[6]), .SP(CS_READY_c_enable_14), 
            .CK(CS_READY_c), .Q(cs_decoded[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i6.GSR = "ENABLED";
    FD1P3AY cs_decoded_i5 (.D(cs_decoded_13__N_752[6]), .SP(CS_READY_c_enable_15), 
            .CK(CS_READY_c), .Q(cs_decoded[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i5.GSR = "ENABLED";
    FD1P3AY cs_decoded_i4 (.D(cs_decoded_13__N_752[6]), .SP(CS_READY_c_enable_16), 
            .CK(CS_READY_c), .Q(cs_decoded[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=213, LSE_RLINE=221 */ ;   // c:/s_links/sources/cs_decoder.v(31[11] 75[5])
    defparam cs_decoded_i4.GSR = "ENABLED";
    LUT4 i2_1_lut (.A(cs_c_4), .Z(FLASH_CS_N_768)) /* synthesis lut_function=(!(A)) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i2_1_lut.init = 16'h5555;
    LUT4 cs_c_0_bdd_4_lut (.A(cs_c_2), .B(cs_c_1), .C(cs_c_4), .D(cs_c_3), 
         .Z(n28852)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;
    defparam cs_c_0_bdd_4_lut.init = 16'h8001;
    LUT4 i1_4_lut (.A(cs_c_1), .B(n29131), .C(n29274), .D(cs_c_2), .Z(CS_READY_c_enable_7)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_4_lut.init = 16'hc8c0;
    LUT4 i22417_4_lut (.A(n29131), .B(n29236), .C(n29274), .D(cs_c_2), 
         .Z(CS_READY_c_enable_9)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i22417_4_lut.init = 16'ha2a0;
    LUT4 i1_4_lut_adj_952 (.A(cs_c_1), .B(n29131), .C(n29274), .D(cs_c_0), 
         .Z(CS_READY_c_enable_10)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i1_4_lut_adj_952.init = 16'hc8c0;
    LUT4 i22419_4_lut (.A(n29131), .B(n27728), .C(n29274), .D(cs_c_1), 
         .Z(CS_READY_c_enable_11)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i22419_4_lut.init = 16'ha2a0;
    LUT4 i22569_2_lut (.A(cs_c_2), .B(cs_c_0), .Z(n27728)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i22569_2_lut.init = 16'h6666;
    LUT4 i22418_4_lut (.A(n29131), .B(n27736), .C(n29274), .D(cs_c_0), 
         .Z(CS_READY_c_enable_12)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i22418_4_lut.init = 16'ha2a0;
    LUT4 i22577_2_lut (.A(cs_c_1), .B(cs_c_2), .Z(n27736)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i22577_2_lut.init = 16'h6666;
    LUT4 i2_4_lut_adj_953 (.A(cs_c_0), .B(n29133), .C(n29292), .D(n27736), 
         .Z(CS_READY_c_enable_15)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D)))) */ ;
    defparam i2_4_lut_adj_953.init = 16'hc0c4;
    LUT4 i2_4_lut_adj_954 (.A(cs_c_1), .B(n29133), .C(n29292), .D(n27728), 
         .Z(CS_READY_c_enable_16)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D)))) */ ;
    defparam i2_4_lut_adj_954.init = 16'hc0c4;
    LUT4 i22947_4_lut (.A(n29163), .B(cs_c_3), .C(n27352), .D(n29258), 
         .Z(CS_READY_c_enable_4)) /* synthesis lut_function=(!(A+!(B (C)+!B (C+!(D))))) */ ;
    defparam i22947_4_lut.init = 16'h5051;
    LUT4 cs_4__I_0_16_Mux_2_i31_4_lut (.A(cs_c_3), .B(n29188), .C(cs_c_4), 
         .D(cs_c_1), .Z(cs_decoded_13__N_752[2])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+(D))+!B !(C+!(D))))) */ ;   // c:/s_links/sources/cs_decoder.v(32[5] 74[10])
    defparam cs_4__I_0_16_Mux_2_i31_4_lut.init = 16'h3a3f;
    LUT4 i1_4_lut_then_4_lut (.A(cs_c_1), .B(cs_c_3), .C(cs_c_2), .D(cs_c_0), 
         .Z(n29331)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_4_lut_then_4_lut.init = 16'h4000;
    LUT4 i22943_4_lut (.A(n29163), .B(cs_c_0), .C(n27352), .D(n27513), 
         .Z(CS_READY_c_enable_6)) /* synthesis lut_function=(!(A+!(B (C)+!B (C+!(D))))) */ ;
    defparam i22943_4_lut.init = 16'h5051;
    LUT4 cs_4__I_0_16_Mux_3_i31_4_lut (.A(cs_c_3), .B(n29188), .C(cs_c_4), 
         .D(cs_c_2), .Z(cs_decoded_13__N_752[3])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+(D))+!B !(C+!(D))))) */ ;   // c:/s_links/sources/cs_decoder.v(32[5] 74[10])
    defparam cs_4__I_0_16_Mux_3_i31_4_lut.init = 16'h3a3f;
    LUT4 i22363_2_lut (.A(cs_c_3), .B(cs_c_1), .Z(n27513)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22363_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_else_4_lut (.A(cs_c_1), .B(cs_c_3), .C(cs_c_2), .D(cs_c_0), 
         .Z(n29330)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/s_links/sources/mcm_top.v(19[37:39])
    defparam i1_4_lut_else_4_lut.init = 16'h0001;
    LUT4 i22945_4_lut_4_lut (.A(n29163), .B(n29292), .C(n33), .D(n29159), 
         .Z(CS_READY_c_enable_5)) /* synthesis lut_function=(!(A+!(B (D)+!B (C (D))))) */ ;
    defparam i22945_4_lut_4_lut.init = 16'h5400;
    LUT4 i1_3_lut_4_lut_adj_955 (.A(n29163), .B(n13889), .C(n29274), .D(n29273), 
         .Z(CS_READY_c_enable_8)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_955.init = 16'h4440;
    LUT4 i108_3_lut_4_lut (.A(n29163), .B(n13889), .C(n29274), .D(n71), 
         .Z(CS_READY_c_enable_13)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i108_3_lut_4_lut.init = 16'h4440;
    
endmodule
//
// Verilog Description of module \intrpt_ctrl(DEV_ID=1) 
//

module \intrpt_ctrl(DEV_ID=1)  (clk, n29239, \spi_data_out_r_39__N_2643[0] , 
            \pin_intrpt[3] , intrpt_out_c_1, intrpt_out_N_2706, n29757, 
            clear_intrpt, clear_intrpt_N_2710, \spi_data_out_r_39__N_2643[2] , 
            \pin_intrpt[5] , \spi_data_out_r_39__N_2643[1] , \pin_intrpt[4] ) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input n29239;
    output \spi_data_out_r_39__N_2643[0] ;
    input \pin_intrpt[3] ;
    output intrpt_out_c_1;
    input intrpt_out_N_2706;
    input n29757;
    output clear_intrpt;
    input clear_intrpt_N_2710;
    output \spi_data_out_r_39__N_2643[2] ;
    input \pin_intrpt[5] ;
    output \spi_data_out_r_39__N_2643[1] ;
    input \pin_intrpt[4] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire \pin_intrpt[5]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[5] */ ;   // c:/s_links/sources/mcm_top.v(102[46:56])
    wire [2:0]intrpt_in_dly;   // c:/s_links/sources/intrpt_ctrl.v(39[36:49])
    wire [2:0]intrpt_in_reg;   // c:/s_links/sources/intrpt_ctrl.v(38[35:48])
    
    wire assert_intrpt, intrpt_all_edges, n4;
    
    FD1S3IX intrpt_in_dly__i0 (.D(intrpt_in_reg[0]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\pin_intrpt[3] ), .CK(clk), .Q(\spi_data_out_r_39__N_2643[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i0 (.D(\pin_intrpt[3] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i0.GSR = "DISABLED";
    FD1P3IX intrpt_out_359 (.D(n29757), .SP(assert_intrpt), .CD(intrpt_out_N_2706), 
            .CK(clk), .Q(intrpt_out_c_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(92[8] 99[4])
    defparam intrpt_out_359.GSR = "DISABLED";
    FD1S3IX clear_intrpt_317 (.D(clear_intrpt_N_2710), .CK(clk), .CD(n29239), 
            .Q(clear_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam clear_intrpt_317.GSR = "DISABLED";
    FD1S3IX assert_intrpt_316 (.D(intrpt_all_edges), .CK(clk), .CD(n29239), 
            .Q(assert_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(63[8] 73[4])
    defparam assert_intrpt_316.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\pin_intrpt[5] ), .CK(clk), .Q(\spi_data_out_r_39__N_2643[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\pin_intrpt[4] ), .CK(clk), .Q(\spi_data_out_r_39__N_2643[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i2 (.D(intrpt_in_reg[2]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i1 (.D(intrpt_in_reg[1]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i1 (.D(\pin_intrpt[4] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i2 (.D(\pin_intrpt[5] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i2.GSR = "DISABLED";
    LUT4 i2_3_lut (.A(intrpt_in_dly[0]), .B(n4), .C(intrpt_in_reg[0]), 
         .Z(intrpt_all_edges)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i2_3_lut.init = 16'hdede;
    LUT4 i1_4_lut (.A(intrpt_in_dly[1]), .B(intrpt_in_dly[2]), .C(intrpt_in_reg[1]), 
         .D(intrpt_in_reg[2]), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i1_4_lut.init = 16'h7bde;
    
endmodule
//
// Verilog Description of module intrpt_ctrl
//

module intrpt_ctrl (\spi_data_out_r_39__N_2572[0] , clk, \pin_intrpt[0] , 
            n29239, intrpt_out_c_0, intrpt_out_N_2635, n29757, clear_intrpt, 
            clear_intrpt_N_2639, n29212, \spi_cmd[2] , n29126, \spi_addr[0] , 
            clear_intrpt_N_2781, clear_intrpt_N_2852, n29178, n29141, 
            \spi_cmd[1] , clear_intrpt_N_2923, clear_intrpt_N_2994, \spi_data_out_r_39__N_2572[2] , 
            \mode[2]_derived_32 , \spi_data_out_r_39__N_2572[1] , \pin_intrpt[1] , 
            n29761, \spi_addr[1] , n29310, \spi_addr[2] , n13413) /* synthesis syn_module_defined=1 */ ;
    output \spi_data_out_r_39__N_2572[0] ;
    input clk;
    input \pin_intrpt[0] ;
    input n29239;
    output intrpt_out_c_0;
    input intrpt_out_N_2635;
    input n29757;
    output clear_intrpt;
    input clear_intrpt_N_2639;
    output n29212;
    input \spi_cmd[2] ;
    input n29126;
    input \spi_addr[0] ;
    output clear_intrpt_N_2781;
    output clear_intrpt_N_2852;
    input n29178;
    input n29141;
    input \spi_cmd[1] ;
    output clear_intrpt_N_2923;
    output clear_intrpt_N_2994;
    output \spi_data_out_r_39__N_2572[2] ;
    input \mode[2]_derived_32 ;
    output \spi_data_out_r_39__N_2572[1] ;
    input \pin_intrpt[1] ;
    input n29761;
    input \spi_addr[1] ;
    output n29310;
    input \spi_addr[2] ;
    output n13413;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire \mode[2]_derived_32  /* synthesis is_clock=1, SET_AS_NETWORK=\stepper_ins[0].u_stepper/mode[2]_derived_32 */ ;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    wire [2:0]intrpt_in_reg;   // c:/s_links/sources/intrpt_ctrl.v(38[35:48])
    wire [2:0]intrpt_in_dly;   // c:/s_links/sources/intrpt_ctrl.v(39[36:49])
    
    wire assert_intrpt, intrpt_all_edges, n4;
    
    FD1S3AX spi_data_out_r_i1 (.D(\pin_intrpt[0] ), .CK(clk), .Q(\spi_data_out_r_39__N_2572[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i0 (.D(\pin_intrpt[0] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i0.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i0 (.D(intrpt_in_reg[0]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i0.GSR = "DISABLED";
    FD1P3IX intrpt_out_359 (.D(n29757), .SP(assert_intrpt), .CD(intrpt_out_N_2635), 
            .CK(clk), .Q(intrpt_out_c_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(92[8] 99[4])
    defparam intrpt_out_359.GSR = "DISABLED";
    FD1S3IX clear_intrpt_317 (.D(clear_intrpt_N_2639), .CK(clk), .CD(n29239), 
            .Q(clear_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam clear_intrpt_317.GSR = "DISABLED";
    FD1S3IX assert_intrpt_316 (.D(intrpt_all_edges), .CK(clk), .CD(n29239), 
            .Q(assert_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(63[8] 73[4])
    defparam assert_intrpt_316.GSR = "DISABLED";
    LUT4 i22921_2_lut_3_lut_4_lut_4_lut (.A(n29212), .B(\spi_cmd[2] ), .C(n29126), 
         .D(\spi_addr[0] ), .Z(clear_intrpt_N_2781)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(82[15:43])
    defparam i22921_2_lut_3_lut_4_lut_4_lut.init = 16'h0001;
    LUT4 i22918_2_lut_3_lut_4_lut_4_lut (.A(n29212), .B(\spi_cmd[2] ), .C(n29126), 
         .D(\spi_addr[0] ), .Z(clear_intrpt_N_2852)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(82[15:43])
    defparam i22918_2_lut_3_lut_4_lut_4_lut.init = 16'h0100;
    LUT4 i22909_2_lut_3_lut_4_lut_4_lut (.A(n29178), .B(\spi_addr[0] ), 
         .C(n29141), .D(\spi_cmd[1] ), .Z(clear_intrpt_N_2923)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(82[15:43])
    defparam i22909_2_lut_3_lut_4_lut_4_lut.init = 16'h0100;
    LUT4 i22906_2_lut_3_lut_4_lut_4_lut (.A(n29178), .B(\spi_addr[0] ), 
         .C(n29141), .D(\spi_cmd[1] ), .Z(clear_intrpt_N_2994)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(82[15:43])
    defparam i22906_2_lut_3_lut_4_lut_4_lut.init = 16'h0400;
    FD1S3AX spi_data_out_r_i3 (.D(\mode[2]_derived_32 ), .CK(clk), .Q(\spi_data_out_r_39__N_2572[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\pin_intrpt[1] ), .CK(clk), .Q(\spi_data_out_r_39__N_2572[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i1 (.D(\pin_intrpt[1] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i2 (.D(\mode[2]_derived_32 ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i1 (.D(intrpt_in_reg[1]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i2 (.D(intrpt_in_reg[2]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i2.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_582 (.A(n29761), .B(\spi_addr[1] ), .Z(n29310)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/intrpt_ctrl.v(82[15:43])
    defparam i1_2_lut_rep_582.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_484_3_lut (.A(n29761), .B(\spi_addr[1] ), .C(\spi_addr[2] ), 
         .Z(n29212)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/s_links/sources/intrpt_ctrl.v(82[15:43])
    defparam i1_2_lut_rep_484_3_lut.init = 16'hfbfb;
    LUT4 i2_3_lut (.A(intrpt_in_dly[0]), .B(n4), .C(intrpt_in_reg[0]), 
         .Z(intrpt_all_edges)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i2_3_lut.init = 16'hdede;
    LUT4 i1_4_lut (.A(intrpt_in_dly[1]), .B(intrpt_in_dly[2]), .C(intrpt_in_reg[1]), 
         .D(intrpt_in_reg[2]), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i1_4_lut.init = 16'h7bde;
    LUT4 i2_3_lut_adj_945 (.A(\spi_addr[1] ), .B(n29761), .C(\spi_addr[2] ), 
         .Z(n13413)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/s_links/sources/intrpt_ctrl.v(82[15:43])
    defparam i2_3_lut_adj_945.init = 16'hf7f7;
    
endmodule
//
// Verilog Description of module quad_decoder
//

module quad_decoder (n29099, n25293, quad_buffer, quad_count, \spi_data_out_r_39__N_2483[9] , 
            \spi_data_out_r_39__N_2483[8] , clk_1MHz, clk_1MHz_enable_340, 
            \spi_data_out_r_39__N_934[0] , clk, \quad_b[0] , \mode[2]_derived_32 , 
            \spi_data_out_r_39__N_2483[7] , \spi_data_out_r_39__N_2483[6] , 
            \spi_data_out_r_39__N_2483[5] , \spi_data_out_r_39__N_2483[4] , 
            \spi_data_out_r_39__N_2483[3] , \spi_data_out_r_39__N_2483[2] , 
            n13413, quad_buffer_adj_528, quad_count_adj_529, \spi_data_out_r_39__N_1547[29] , 
            \spi_data_out_r_39__N_2483[1] , n29239, \spi_addr[1] , n29761, 
            \spi_addr[2] , n13506, n13511, \spi_data_out_r_39__N_1547[28] , 
            clk_enable_433, \spi_data_r[0] , quad_homing, clk_enable_436, 
            n29762, n29098, quad_buffer_adj_530, quad_count_adj_531, 
            \spi_data_out_r_39__N_2249[0] , \spi_data_out_r_39__N_2249[31] , 
            \spi_data_out_r_39__N_2249[30] , \spi_data_out_r_39__N_2249[29] , 
            \spi_data_out_r_39__N_2249[28] , \spi_data_out_r_39__N_2249[27] , 
            \spi_data_out_r_39__N_2249[26] , \spi_data_out_r_39__N_2249[25] , 
            \spi_data_out_r_39__N_2249[24] , \spi_data_out_r_39__N_2249[23] , 
            \spi_data_out_r_39__N_2249[22] , \spi_data_out_r_39__N_1547[27] , 
            \spi_data_out_r_39__N_2249[21] , \spi_data_out_r_39__N_2249[20] , 
            quad_buffer_adj_532, quad_count_adj_533, \spi_data_out_r_39__N_2015[27] , 
            \spi_data_out_r_39__N_2015[26] , \spi_data_out_r_39__N_2015[25] , 
            \spi_data_out_r_39__N_2015[24] , \spi_data_out_r_39__N_2015[23] , 
            \spi_data_out_r_39__N_2249[19] , \spi_data_out_r_39__N_2249[18] , 
            \spi_data_out_r_39__N_1547[26] , \spi_data_out_r_39__N_1547[25] , 
            \spi_data_out_r_39__N_2249[17] , \spi_data_out_r_39__N_2015[22] , 
            \spi_data_out_r_39__N_2249[16] , \spi_data_out_r_39__N_2249[15] , 
            \spi_data_out_r_39__N_1547[24] , \spi_data_out_r_39__N_2249[14] , 
            \spi_data_out_r_39__N_2015[21] , \spi_data_out_r_39__N_2015[20] , 
            \spi_data_out_r_39__N_2249[13] , \spi_data_out_r_39__N_2015[19] , 
            \spi_data_out_r_39__N_2015[18] , \spi_data_out_r_39__N_2015[17] , 
            \spi_data_out_r_39__N_2249[12] , \spi_data_out_r_39__N_2015[16] , 
            \spi_data_out_r_39__N_2015[15] , \spi_data_out_r_39__N_2015[14] , 
            \spi_data_out_r_39__N_2015[13] , \spi_data_out_r_39__N_2249[11] , 
            \spi_data_out_r_39__N_2249[10] , \spi_data_out_r_39__N_2249[9] , 
            spi_data_out_r_39__N_974, spi_data_out_r_39__N_1162, \spi_data_out_r_39__N_2249[8] , 
            quad_set_complete, quad_set_valid, \spi_data_out_r_39__N_2015[12] , 
            \spi_data_out_r_39__N_2015[11] , \spi_data_out_r_39__N_2249[7] , 
            \spi_data_out_r_39__N_2249[6] , \spi_data_out_r_39__N_2249[5] , 
            \spi_data_out_r_39__N_2249[4] , \spi_data_out_r_39__N_1547[23] , 
            \spi_data_out_r_39__N_2015[10] , \spi_data_out_r_39__N_2015[9] , 
            \spi_data_out_r_39__N_2249[3] , \spi_data_out_r_39__N_2015[8] , 
            \spi_data_out_r_39__N_2015[7] , \spi_data_out_r_39__N_2015[6] , 
            \spi_data_out_r_39__N_2015[5] , \spi_data_out_r_39__N_1547[22] , 
            \spi_data_out_r_39__N_2249[2] , \spi_data_out_r_39__N_1547[21] , 
            \spi_data_out_r_39__N_2015[4] , \spi_data_out_r_39__N_2015[3] , 
            \spi_data_out_r_39__N_1547[20] , \spi_data_out_r_39__N_2249[1] , 
            \spi_data_out_r_39__N_2015[2] , \spi_data_out_r_39__N_2015[1] , 
            quad_buffer_adj_534, quad_count_adj_535, \spi_data_out_r_39__N_1781[0] , 
            \spi_data_out_r_39__N_1547[19] , \spi_data_out_r_39__N_1781[31] , 
            \spi_data_out_r_39__N_1781[30] , \spi_data_out_r_39__N_1781[29] , 
            \spi_data_out_r_39__N_1781[28] , \spi_data_out_r_39__N_1781[27] , 
            n29260, pin_io_out_4, n108, n79, \spi_data_out_r_39__N_1781[26] , 
            \spi_data_out_r_39__N_1547[18] , \spi_data_out_r_39__N_1547[17] , 
            \spi_data_out_r_39__N_1781[25] , \spi_data_out_r_39__N_1781[24] , 
            \spi_data_out_r_39__N_1781[23] , \spi_data_out_r_39__N_1547[16] , 
            \spi_data_out_r_39__N_1781[22] , \spi_data_out_r_39__N_1781[21] , 
            \spi_data_out_r_39__N_1781[20] , \spi_data_out_r_39__N_1781[19] , 
            \spi_data_out_r_39__N_1781[18] , \spi_data_out_r_39__N_1547[15] , 
            \spi_data_out_r_39__N_1547[14] , \spi_data_out_r_39__N_1781[17] , 
            \spi_data_out_r_39__N_1781[16] , \spi_data_out_r_39__N_1781[15] , 
            \spi_data_out_r_39__N_1781[14] , \spi_data_out_r_39__N_1781[13] , 
            \spi_data_out_r_39__N_1781[12] , \spi_data_out_r_39__N_1781[11] , 
            \spi_data_out_r_39__N_1547[13] , \spi_data_out_r_39__N_1781[10] , 
            \spi_data_out_r_39__N_1781[9] , \spi_data_out_r_39__N_1781[8] , 
            \spi_data_out_r_39__N_1781[7] , \spi_data_out_r_39__N_1781[6] , 
            \spi_data_out_r_39__N_1781[5] , n27256, n29078, n27338, 
            n29213, clk_enable_199, \spi_data_out_r_39__N_1781[4] , \spi_data_out_r_39__N_1781[3] , 
            \spi_data_out_r_39__N_1781[2] , \spi_data_out_r_39__N_1781[1] , 
            \spi_data_out_r_39__N_2483[0] , \spi_data_out_r_39__N_2483[31] , 
            \spi_data_out_r_39__N_2483[30] , \spi_data_out_r_39__N_2483[29] , 
            \spi_data_out_r_39__N_2483[28] , \spi_data_out_r_39__N_1547[0] , 
            \spi_data_out_r_39__N_2483[27] , \spi_data_out_r_39__N_2483[26] , 
            resetn_c, GND_net, \spi_data_out_r_39__N_2483[25] , \spi_data_out_r_39__N_2483[24] , 
            \spi_data_out_r_39__N_2483[23] , \spi_data_out_r_39__N_2483[22] , 
            \spi_data_out_r_39__N_2483[21] , \spi_data_out_r_39__N_2483[20] , 
            \spi_data_out_r_39__N_2483[19] , \spi_data_out_r_39__N_2483[18] , 
            \spi_data_out_r_39__N_2483[17] , \spi_data_out_r_39__N_1547[12] , 
            \spi_data_out_r_39__N_2483[16] , \spi_data_out_r_39__N_1547[31] , 
            \spi_data_out_r_39__N_2483[15] , \spi_data_out_r_39__N_1547[30] , 
            \spi_data_out_r_39__N_2483[14] , \spi_data_out_r_39__N_1547[11] , 
            \spi_data_out_r_39__N_1547[10] , \spi_data_out_r_39__N_2483[13] , 
            \spi_data_out_r_39__N_1547[9] , \spi_data_out_r_39__N_2483[12] , 
            \spi_data_out_r_39__N_2483[11] , \spi_data_out_r_39__N_2483[10] , 
            \spi_data_out_r_39__N_1547[8] , \quad_a[0] , \spi_data_out_r_39__N_934[31] , 
            \spi_data_out_r_39__N_934[30] , \spi_data_out_r_39__N_934[29] , 
            \spi_data_out_r_39__N_1547[7] , \spi_data_out_r_39__N_934[28] , 
            \spi_data_out_r_39__N_934[27] , \spi_data_out_r_39__N_934[26] , 
            \spi_data_out_r_39__N_934[25] , \spi_data_out_r_39__N_934[24] , 
            \spi_data_out_r_39__N_934[23] , \spi_data_out_r_39__N_934[22] , 
            \spi_data_out_r_39__N_934[21] , \spi_data_out_r_39__N_934[20] , 
            \spi_data_out_r_39__N_934[19] , \spi_data_out_r_39__N_934[18] , 
            \spi_data_out_r_39__N_934[17] , \spi_data_out_r_39__N_934[16] , 
            \spi_data_out_r_39__N_934[15] , \spi_data_out_r_39__N_934[14] , 
            \spi_data_out_r_39__N_934[13] , \spi_data_out_r_39__N_934[12] , 
            \spi_data_out_r_39__N_934[11] , \spi_data_out_r_39__N_934[10] , 
            \spi_data_out_r_39__N_934[9] , \spi_data_out_r_39__N_934[8] , 
            \spi_data_out_r_39__N_934[7] , \spi_data_out_r_39__N_934[6] , 
            \spi_data_out_r_39__N_934[5] , \spi_data_out_r_39__N_934[4] , 
            \spi_data_out_r_39__N_934[3] , \spi_data_out_r_39__N_934[2] , 
            \spi_data_out_r_39__N_934[1] , \spi_data_out_r_39__N_1547[6] , 
            \spi_data_out_r_39__N_1547[5] , \spi_data_out_r_39__N_1547[4] , 
            \spi_data_out_r_39__N_1547[3] , \spi_data_out_r_39__N_1547[2] , 
            \spi_data_out_r_39__N_1547[1] , quad_buffer_adj_536, quad_count_adj_537, 
            \spi_data_out_r_39__N_1313[0] , \spi_data_out_r_39__N_1313[31] , 
            \spi_cmd[2] , n29117, n29310, clear_intrpt_N_3065, \spi_data_out_r_39__N_1313[30] , 
            \spi_data_out_r_39__N_1313[29] , \spi_data_out_r_39__N_1313[28] , 
            \spi_data_out_r_39__N_1313[27] , \spi_data_r[1] , \spi_data_r[2] , 
            \spi_data_r[3] , \spi_data_r[4] , \spi_data_r[5] , \spi_data_r[6] , 
            \spi_data_r[7] , \spi_data_r[8] , \spi_data_r[9] , \spi_data_r[10] , 
            \spi_data_r[11] , \spi_data_r[12] , \spi_data_r[13] , \spi_data_r[14] , 
            \spi_data_r[15] , \spi_data_r[16] , \spi_data_r[17] , \spi_data_r[18] , 
            \spi_data_r[19] , \spi_data_r[20] , \spi_data_r[21] , \spi_data_r[22] , 
            \spi_data_r[23] , \spi_data_r[24] , \spi_data_r[25] , \spi_data_r[26] , 
            \spi_data_r[27] , \spi_data_r[28] , \spi_data_r[29] , \spi_data_r[30] , 
            \spi_data_r[31] , clk_enable_501, n29085, \spi_data_out_r_39__N_1313[26] , 
            \spi_data_out_r_39__N_1313[25] , \spi_data_out_r_39__N_1313[24] , 
            n3, n26, \spi_data_out_r_39__N_1313[23] , \spi_data_out_r_39__N_1313[22] , 
            \spi_data_out_r_39__N_1313[21] , \spi_data_out_r_39__N_1313[20] , 
            \spi_data_out_r_39__N_1313[19] , \spi_data_out_r_39__N_1313[18] , 
            \spi_data_out_r_39__N_1313[17] , n20819, \spi_data_out_r_39__N_1313[16] , 
            \spi_data_out_r_39__N_1313[15] , \spi_data_out_r_39__N_1313[14] , 
            n31, \spi_data_out_r_39__N_1313[13] , \spi_data_out_r_39__N_1313[12] , 
            \spi_data_out_r_39__N_1313[11] , \spi_data_out_r_39__N_1313[10] , 
            \spi_data_out_r_39__N_1313[9] , \spi_data_out_r_39__N_1313[8] , 
            \spi_data_out_r_39__N_1313[7] , \spi_data_out_r_39__N_1313[6] , 
            \spi_data_out_r_39__N_1313[5] , \spi_data_out_r_39__N_1313[4] , 
            \spi_data_out_r_39__N_1313[3] , \spi_data_out_r_39__N_1313[2] , 
            \spi_data_out_r_39__N_1313[1] , \spi_data_out_r_39__N_2015[0] , 
            \spi_data_out_r_39__N_2015[31] , \spi_data_out_r_39__N_2015[30] , 
            \spi_data_out_r_39__N_2015[29] , n29326, \spi_data_out_r_39__N_2015[28] ) /* synthesis syn_module_defined=1 */ ;
    input n29099;
    output n25293;
    input [31:0]quad_buffer;
    input [31:0]quad_count;
    output \spi_data_out_r_39__N_2483[9] ;
    output \spi_data_out_r_39__N_2483[8] ;
    input clk_1MHz;
    input clk_1MHz_enable_340;
    output \spi_data_out_r_39__N_934[0] ;
    input clk;
    input \quad_b[0] ;
    input \mode[2]_derived_32 ;
    output \spi_data_out_r_39__N_2483[7] ;
    output \spi_data_out_r_39__N_2483[6] ;
    output \spi_data_out_r_39__N_2483[5] ;
    output \spi_data_out_r_39__N_2483[4] ;
    output \spi_data_out_r_39__N_2483[3] ;
    output \spi_data_out_r_39__N_2483[2] ;
    input n13413;
    input [31:0]quad_buffer_adj_528;
    input [31:0]quad_count_adj_529;
    output \spi_data_out_r_39__N_1547[29] ;
    output \spi_data_out_r_39__N_2483[1] ;
    input n29239;
    input \spi_addr[1] ;
    input n29761;
    input \spi_addr[2] ;
    output n13506;
    output n13511;
    output \spi_data_out_r_39__N_1547[28] ;
    input clk_enable_433;
    input \spi_data_r[0] ;
    output [1:0]quad_homing;
    input clk_enable_436;
    input n29762;
    input n29098;
    input [31:0]quad_buffer_adj_530;
    input [31:0]quad_count_adj_531;
    output \spi_data_out_r_39__N_2249[0] ;
    output \spi_data_out_r_39__N_2249[31] ;
    output \spi_data_out_r_39__N_2249[30] ;
    output \spi_data_out_r_39__N_2249[29] ;
    output \spi_data_out_r_39__N_2249[28] ;
    output \spi_data_out_r_39__N_2249[27] ;
    output \spi_data_out_r_39__N_2249[26] ;
    output \spi_data_out_r_39__N_2249[25] ;
    output \spi_data_out_r_39__N_2249[24] ;
    output \spi_data_out_r_39__N_2249[23] ;
    output \spi_data_out_r_39__N_2249[22] ;
    output \spi_data_out_r_39__N_1547[27] ;
    output \spi_data_out_r_39__N_2249[21] ;
    output \spi_data_out_r_39__N_2249[20] ;
    input [31:0]quad_buffer_adj_532;
    input [31:0]quad_count_adj_533;
    output \spi_data_out_r_39__N_2015[27] ;
    output \spi_data_out_r_39__N_2015[26] ;
    output \spi_data_out_r_39__N_2015[25] ;
    output \spi_data_out_r_39__N_2015[24] ;
    output \spi_data_out_r_39__N_2015[23] ;
    output \spi_data_out_r_39__N_2249[19] ;
    output \spi_data_out_r_39__N_2249[18] ;
    output \spi_data_out_r_39__N_1547[26] ;
    output \spi_data_out_r_39__N_1547[25] ;
    output \spi_data_out_r_39__N_2249[17] ;
    output \spi_data_out_r_39__N_2015[22] ;
    output \spi_data_out_r_39__N_2249[16] ;
    output \spi_data_out_r_39__N_2249[15] ;
    output \spi_data_out_r_39__N_1547[24] ;
    output \spi_data_out_r_39__N_2249[14] ;
    output \spi_data_out_r_39__N_2015[21] ;
    output \spi_data_out_r_39__N_2015[20] ;
    output \spi_data_out_r_39__N_2249[13] ;
    output \spi_data_out_r_39__N_2015[19] ;
    output \spi_data_out_r_39__N_2015[18] ;
    output \spi_data_out_r_39__N_2015[17] ;
    output \spi_data_out_r_39__N_2249[12] ;
    output \spi_data_out_r_39__N_2015[16] ;
    output \spi_data_out_r_39__N_2015[15] ;
    output \spi_data_out_r_39__N_2015[14] ;
    output \spi_data_out_r_39__N_2015[13] ;
    output \spi_data_out_r_39__N_2249[11] ;
    output \spi_data_out_r_39__N_2249[10] ;
    output \spi_data_out_r_39__N_2249[9] ;
    output spi_data_out_r_39__N_974;
    input spi_data_out_r_39__N_1162;
    output \spi_data_out_r_39__N_2249[8] ;
    output quad_set_complete;
    output quad_set_valid;
    output \spi_data_out_r_39__N_2015[12] ;
    output \spi_data_out_r_39__N_2015[11] ;
    output \spi_data_out_r_39__N_2249[7] ;
    output \spi_data_out_r_39__N_2249[6] ;
    output \spi_data_out_r_39__N_2249[5] ;
    output \spi_data_out_r_39__N_2249[4] ;
    output \spi_data_out_r_39__N_1547[23] ;
    output \spi_data_out_r_39__N_2015[10] ;
    output \spi_data_out_r_39__N_2015[9] ;
    output \spi_data_out_r_39__N_2249[3] ;
    output \spi_data_out_r_39__N_2015[8] ;
    output \spi_data_out_r_39__N_2015[7] ;
    output \spi_data_out_r_39__N_2015[6] ;
    output \spi_data_out_r_39__N_2015[5] ;
    output \spi_data_out_r_39__N_1547[22] ;
    output \spi_data_out_r_39__N_2249[2] ;
    output \spi_data_out_r_39__N_1547[21] ;
    output \spi_data_out_r_39__N_2015[4] ;
    output \spi_data_out_r_39__N_2015[3] ;
    output \spi_data_out_r_39__N_1547[20] ;
    output \spi_data_out_r_39__N_2249[1] ;
    output \spi_data_out_r_39__N_2015[2] ;
    output \spi_data_out_r_39__N_2015[1] ;
    input [31:0]quad_buffer_adj_534;
    input [31:0]quad_count_adj_535;
    output \spi_data_out_r_39__N_1781[0] ;
    output \spi_data_out_r_39__N_1547[19] ;
    output \spi_data_out_r_39__N_1781[31] ;
    output \spi_data_out_r_39__N_1781[30] ;
    output \spi_data_out_r_39__N_1781[29] ;
    output \spi_data_out_r_39__N_1781[28] ;
    output \spi_data_out_r_39__N_1781[27] ;
    input n29260;
    input pin_io_out_4;
    output n108;
    output n79;
    output \spi_data_out_r_39__N_1781[26] ;
    output \spi_data_out_r_39__N_1547[18] ;
    output \spi_data_out_r_39__N_1547[17] ;
    output \spi_data_out_r_39__N_1781[25] ;
    output \spi_data_out_r_39__N_1781[24] ;
    output \spi_data_out_r_39__N_1781[23] ;
    output \spi_data_out_r_39__N_1547[16] ;
    output \spi_data_out_r_39__N_1781[22] ;
    output \spi_data_out_r_39__N_1781[21] ;
    output \spi_data_out_r_39__N_1781[20] ;
    output \spi_data_out_r_39__N_1781[19] ;
    output \spi_data_out_r_39__N_1781[18] ;
    output \spi_data_out_r_39__N_1547[15] ;
    output \spi_data_out_r_39__N_1547[14] ;
    output \spi_data_out_r_39__N_1781[17] ;
    output \spi_data_out_r_39__N_1781[16] ;
    output \spi_data_out_r_39__N_1781[15] ;
    output \spi_data_out_r_39__N_1781[14] ;
    output \spi_data_out_r_39__N_1781[13] ;
    output \spi_data_out_r_39__N_1781[12] ;
    output \spi_data_out_r_39__N_1781[11] ;
    output \spi_data_out_r_39__N_1547[13] ;
    output \spi_data_out_r_39__N_1781[10] ;
    output \spi_data_out_r_39__N_1781[9] ;
    output \spi_data_out_r_39__N_1781[8] ;
    output \spi_data_out_r_39__N_1781[7] ;
    output \spi_data_out_r_39__N_1781[6] ;
    output \spi_data_out_r_39__N_1781[5] ;
    input n27256;
    input n29078;
    input n27338;
    input n29213;
    output clk_enable_199;
    output \spi_data_out_r_39__N_1781[4] ;
    output \spi_data_out_r_39__N_1781[3] ;
    output \spi_data_out_r_39__N_1781[2] ;
    output \spi_data_out_r_39__N_1781[1] ;
    output \spi_data_out_r_39__N_2483[0] ;
    output \spi_data_out_r_39__N_2483[31] ;
    output \spi_data_out_r_39__N_2483[30] ;
    output \spi_data_out_r_39__N_2483[29] ;
    output \spi_data_out_r_39__N_2483[28] ;
    output \spi_data_out_r_39__N_1547[0] ;
    output \spi_data_out_r_39__N_2483[27] ;
    output \spi_data_out_r_39__N_2483[26] ;
    input resetn_c;
    input GND_net;
    output \spi_data_out_r_39__N_2483[25] ;
    output \spi_data_out_r_39__N_2483[24] ;
    output \spi_data_out_r_39__N_2483[23] ;
    output \spi_data_out_r_39__N_2483[22] ;
    output \spi_data_out_r_39__N_2483[21] ;
    output \spi_data_out_r_39__N_2483[20] ;
    output \spi_data_out_r_39__N_2483[19] ;
    output \spi_data_out_r_39__N_2483[18] ;
    output \spi_data_out_r_39__N_2483[17] ;
    output \spi_data_out_r_39__N_1547[12] ;
    output \spi_data_out_r_39__N_2483[16] ;
    output \spi_data_out_r_39__N_1547[31] ;
    output \spi_data_out_r_39__N_2483[15] ;
    output \spi_data_out_r_39__N_1547[30] ;
    output \spi_data_out_r_39__N_2483[14] ;
    output \spi_data_out_r_39__N_1547[11] ;
    output \spi_data_out_r_39__N_1547[10] ;
    output \spi_data_out_r_39__N_2483[13] ;
    output \spi_data_out_r_39__N_1547[9] ;
    output \spi_data_out_r_39__N_2483[12] ;
    output \spi_data_out_r_39__N_2483[11] ;
    output \spi_data_out_r_39__N_2483[10] ;
    output \spi_data_out_r_39__N_1547[8] ;
    input \quad_a[0] ;
    output \spi_data_out_r_39__N_934[31] ;
    output \spi_data_out_r_39__N_934[30] ;
    output \spi_data_out_r_39__N_934[29] ;
    output \spi_data_out_r_39__N_1547[7] ;
    output \spi_data_out_r_39__N_934[28] ;
    output \spi_data_out_r_39__N_934[27] ;
    output \spi_data_out_r_39__N_934[26] ;
    output \spi_data_out_r_39__N_934[25] ;
    output \spi_data_out_r_39__N_934[24] ;
    output \spi_data_out_r_39__N_934[23] ;
    output \spi_data_out_r_39__N_934[22] ;
    output \spi_data_out_r_39__N_934[21] ;
    output \spi_data_out_r_39__N_934[20] ;
    output \spi_data_out_r_39__N_934[19] ;
    output \spi_data_out_r_39__N_934[18] ;
    output \spi_data_out_r_39__N_934[17] ;
    output \spi_data_out_r_39__N_934[16] ;
    output \spi_data_out_r_39__N_934[15] ;
    output \spi_data_out_r_39__N_934[14] ;
    output \spi_data_out_r_39__N_934[13] ;
    output \spi_data_out_r_39__N_934[12] ;
    output \spi_data_out_r_39__N_934[11] ;
    output \spi_data_out_r_39__N_934[10] ;
    output \spi_data_out_r_39__N_934[9] ;
    output \spi_data_out_r_39__N_934[8] ;
    output \spi_data_out_r_39__N_934[7] ;
    output \spi_data_out_r_39__N_934[6] ;
    output \spi_data_out_r_39__N_934[5] ;
    output \spi_data_out_r_39__N_934[4] ;
    output \spi_data_out_r_39__N_934[3] ;
    output \spi_data_out_r_39__N_934[2] ;
    output \spi_data_out_r_39__N_934[1] ;
    output \spi_data_out_r_39__N_1547[6] ;
    output \spi_data_out_r_39__N_1547[5] ;
    output \spi_data_out_r_39__N_1547[4] ;
    output \spi_data_out_r_39__N_1547[3] ;
    output \spi_data_out_r_39__N_1547[2] ;
    output \spi_data_out_r_39__N_1547[1] ;
    input [31:0]quad_buffer_adj_536;
    input [31:0]quad_count_adj_537;
    output \spi_data_out_r_39__N_1313[0] ;
    output \spi_data_out_r_39__N_1313[31] ;
    input \spi_cmd[2] ;
    input n29117;
    input n29310;
    output clear_intrpt_N_3065;
    output \spi_data_out_r_39__N_1313[30] ;
    output \spi_data_out_r_39__N_1313[29] ;
    output \spi_data_out_r_39__N_1313[28] ;
    output \spi_data_out_r_39__N_1313[27] ;
    input \spi_data_r[1] ;
    input \spi_data_r[2] ;
    input \spi_data_r[3] ;
    input \spi_data_r[4] ;
    input \spi_data_r[5] ;
    input \spi_data_r[6] ;
    input \spi_data_r[7] ;
    input \spi_data_r[8] ;
    input \spi_data_r[9] ;
    input \spi_data_r[10] ;
    input \spi_data_r[11] ;
    input \spi_data_r[12] ;
    input \spi_data_r[13] ;
    input \spi_data_r[14] ;
    input \spi_data_r[15] ;
    input \spi_data_r[16] ;
    input \spi_data_r[17] ;
    input \spi_data_r[18] ;
    input \spi_data_r[19] ;
    input \spi_data_r[20] ;
    input \spi_data_r[21] ;
    input \spi_data_r[22] ;
    input \spi_data_r[23] ;
    input \spi_data_r[24] ;
    input \spi_data_r[25] ;
    input \spi_data_r[26] ;
    input \spi_data_r[27] ;
    input \spi_data_r[28] ;
    input \spi_data_r[29] ;
    input \spi_data_r[30] ;
    input \spi_data_r[31] ;
    input clk_enable_501;
    input n29085;
    output \spi_data_out_r_39__N_1313[26] ;
    output \spi_data_out_r_39__N_1313[25] ;
    output \spi_data_out_r_39__N_1313[24] ;
    input n3;
    input n26;
    output \spi_data_out_r_39__N_1313[23] ;
    output \spi_data_out_r_39__N_1313[22] ;
    output \spi_data_out_r_39__N_1313[21] ;
    output \spi_data_out_r_39__N_1313[20] ;
    output \spi_data_out_r_39__N_1313[19] ;
    output \spi_data_out_r_39__N_1313[18] ;
    output \spi_data_out_r_39__N_1313[17] ;
    output n20819;
    output \spi_data_out_r_39__N_1313[16] ;
    output \spi_data_out_r_39__N_1313[15] ;
    output \spi_data_out_r_39__N_1313[14] ;
    output n31;
    output \spi_data_out_r_39__N_1313[13] ;
    output \spi_data_out_r_39__N_1313[12] ;
    output \spi_data_out_r_39__N_1313[11] ;
    output \spi_data_out_r_39__N_1313[10] ;
    output \spi_data_out_r_39__N_1313[9] ;
    output \spi_data_out_r_39__N_1313[8] ;
    output \spi_data_out_r_39__N_1313[7] ;
    output \spi_data_out_r_39__N_1313[6] ;
    output \spi_data_out_r_39__N_1313[5] ;
    output \spi_data_out_r_39__N_1313[4] ;
    output \spi_data_out_r_39__N_1313[3] ;
    output \spi_data_out_r_39__N_1313[2] ;
    output \spi_data_out_r_39__N_1313[1] ;
    output \spi_data_out_r_39__N_2015[0] ;
    output \spi_data_out_r_39__N_2015[31] ;
    output \spi_data_out_r_39__N_2015[30] ;
    output \spi_data_out_r_39__N_2015[29] ;
    output n29326;
    output \spi_data_out_r_39__N_2015[28] ;
    
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire [1:0]sync /* synthesis ASYNC_REG="TRUE" */ ;   // c:/s_links/sources/quad_decoder.v(106[30:34])
    wire [1:0]AB /* synthesis ASYNC_REG="TRUE" */ ;   // c:/s_links/sources/quad_decoder.v(106[36:38])
    wire \mode[2]_derived_32  /* synthesis is_clock=1, SET_AS_NETWORK=\stepper_ins[0].u_stepper/mode[2]_derived_32 */ ;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    wire [31:0]quad_count_adj_7594;   // c:/s_links/sources/quad_decoder.v(45[29:39])
    
    wire n9438;
    wire [39:0]spi_data_out_r_39__N_1079;
    wire [31:0]quad_buffer_adj_7595;   // c:/s_links/sources/quad_decoder.v(46[29:40])
    wire [3:0]n1331;
    
    wire n51, n41, n29034;
    wire [31:0]quad_set;   // c:/s_links/sources/quad_decoder.v(40[31:39])
    
    wire n29321, n20883, n29259, n4, n29261, n9539, n29322, n9547, 
        n25070;
    wire [31:0]n6496;
    
    wire n25069, n25068, n25067, n25066, n25065, n25064, n25063, 
        n25062, n25061, n25060, n25059, n25058, n25057, n25056, 
        n25055, n29320, n10353, n10355, n10357, n10359, n10361, 
        n10363, n10365, n10367, n10369, n10371, n10373, n10375, 
        n10377, n10379, n10381, n10383, n10385, n10387, n10389, 
        n10391, n10393, n10395, n10397, n10399, n10401, n10403, 
        n10405, n10407, n10409, n10411, n10413;
    
    LUT4 mux_863_i10_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[9]), 
         .D(quad_count[9]), .Z(\spi_data_out_r_39__N_2483[9] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i10_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i9_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[8]), 
         .D(quad_count[8]), .Z(\spi_data_out_r_39__N_2483[8] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i9_3_lut_4_lut.init = 16'hf4b0;
    FD1P3AX quad_count_i0_i0 (.D(n9438), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(spi_data_out_r_39__N_1079[0]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX sync_i0 (.D(\quad_b[0] ), .CK(clk_1MHz), .Q(sync[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam sync_i0.GSR = "DISABLED";
    FD1S3AX AB_i0 (.D(sync[0]), .CK(clk_1MHz), .Q(AB[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam AB_i0.GSR = "DISABLED";
    FD1S3AX quad_buffer_i0 (.D(quad_count_adj_7594[0]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i0.GSR = "DISABLED";
    LUT4 mux_863_i8_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[7]), 
         .D(quad_count[7]), .Z(\spi_data_out_r_39__N_2483[7] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i7_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[6]), 
         .D(quad_count[6]), .Z(\spi_data_out_r_39__N_2483[6] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i6_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[5]), 
         .D(quad_count[5]), .Z(\spi_data_out_r_39__N_2483[5] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i5_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[4]), 
         .D(quad_count[4]), .Z(\spi_data_out_r_39__N_2483[4] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i4_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[3]), 
         .D(quad_count[3]), .Z(\spi_data_out_r_39__N_2483[3] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i3_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[2]), 
         .D(quad_count[2]), .Z(\spi_data_out_r_39__N_2483[2] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i3_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_859_i30_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[29]), 
         .D(quad_count_adj_529[29]), .Z(\spi_data_out_r_39__N_1547[29] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_863_i2_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[1]), 
         .D(quad_count[1]), .Z(\spi_data_out_r_39__N_2483[1] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i30_3_lut_4_lut (.A(AB[1]), .B(AB[0]), .C(n1331[3]), .D(n51), 
         .Z(n41)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam i30_3_lut_4_lut.init = 16'h2f20;
    FD1S3JX state_FSM_i0 (.D(n29034), .CK(clk_1MHz), .PD(n29239), .Q(n1331[0]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i0.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut (.A(\spi_addr[1] ), .B(n29761), .C(\spi_addr[2] ), 
         .Z(n13506)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam i1_2_lut_3_lut.init = 16'hfbfb;
    LUT4 i1_2_lut_3_lut_adj_943 (.A(\spi_addr[1] ), .B(n29761), .C(\spi_addr[2] ), 
         .Z(n13511)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam i1_2_lut_3_lut_adj_943.init = 16'hbfbf;
    LUT4 mux_859_i29_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[28]), 
         .D(quad_count_adj_529[28]), .Z(\spi_data_out_r_39__N_1547[28] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i29_3_lut_4_lut.init = 16'hf1e0;
    FD1P3IX quad_set__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i0.GSR = "DISABLED";
    FD1P3IX quad_homing__i0 (.D(n29762), .SP(clk_enable_436), .CD(n29239), 
            .CK(clk), .Q(quad_homing[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam quad_homing__i0.GSR = "DISABLED";
    LUT4 mux_862_i1_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[0]), 
         .D(quad_count_adj_531[0]), .Z(\spi_data_out_r_39__N_2249[0] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i32_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[31]), 
         .D(quad_count_adj_531[31]), .Z(\spi_data_out_r_39__N_2249[31] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i31_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[30]), 
         .D(quad_count_adj_531[30]), .Z(\spi_data_out_r_39__N_2249[30] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i30_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[29]), 
         .D(quad_count_adj_531[29]), .Z(\spi_data_out_r_39__N_2249[29] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i29_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[28]), 
         .D(quad_count_adj_531[28]), .Z(\spi_data_out_r_39__N_2249[28] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i28_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[27]), 
         .D(quad_count_adj_531[27]), .Z(\spi_data_out_r_39__N_2249[27] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i27_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[26]), 
         .D(quad_count_adj_531[26]), .Z(\spi_data_out_r_39__N_2249[26] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i26_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[25]), 
         .D(quad_count_adj_531[25]), .Z(\spi_data_out_r_39__N_2249[25] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i25_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[24]), 
         .D(quad_count_adj_531[24]), .Z(\spi_data_out_r_39__N_2249[24] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i24_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[23]), 
         .D(quad_count_adj_531[23]), .Z(\spi_data_out_r_39__N_2249[23] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i23_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[22]), 
         .D(quad_count_adj_531[22]), .Z(\spi_data_out_r_39__N_2249[22] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i28_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[27]), 
         .D(quad_count_adj_529[27]), .Z(\spi_data_out_r_39__N_1547[27] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i22_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[21]), 
         .D(quad_count_adj_531[21]), .Z(\spi_data_out_r_39__N_2249[21] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i21_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[20]), 
         .D(quad_count_adj_531[20]), .Z(\spi_data_out_r_39__N_2249[20] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i28_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[27]), 
         .D(quad_count_adj_533[27]), .Z(\spi_data_out_r_39__N_2015[27] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i27_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[26]), 
         .D(quad_count_adj_533[26]), .Z(\spi_data_out_r_39__N_2015[26] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i26_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[25]), 
         .D(quad_count_adj_533[25]), .Z(\spi_data_out_r_39__N_2015[25] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i25_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[24]), 
         .D(quad_count_adj_533[24]), .Z(\spi_data_out_r_39__N_2015[24] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i24_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[23]), 
         .D(quad_count_adj_533[23]), .Z(\spi_data_out_r_39__N_2015[23] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i20_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[19]), 
         .D(quad_count_adj_531[19]), .Z(\spi_data_out_r_39__N_2249[19] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i19_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[18]), 
         .D(quad_count_adj_531[18]), .Z(\spi_data_out_r_39__N_2249[18] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i27_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[26]), 
         .D(quad_count_adj_529[26]), .Z(\spi_data_out_r_39__N_1547[26] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i26_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[25]), 
         .D(quad_count_adj_529[25]), .Z(\spi_data_out_r_39__N_1547[25] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i18_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[17]), 
         .D(quad_count_adj_531[17]), .Z(\spi_data_out_r_39__N_2249[17] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i23_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[22]), 
         .D(quad_count_adj_533[22]), .Z(\spi_data_out_r_39__N_2015[22] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i17_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[16]), 
         .D(quad_count_adj_531[16]), .Z(\spi_data_out_r_39__N_2249[16] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i37_4_lut_then_3_lut (.A(n1331[2]), .B(AB[0]), .C(AB[1]), .Z(n29321)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;
    defparam i37_4_lut_then_3_lut.init = 16'h3838;
    LUT4 mux_862_i16_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[15]), 
         .D(quad_count_adj_531[15]), .Z(\spi_data_out_r_39__N_2249[15] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i15940_4_lut_4_lut_4_lut (.A(AB[0]), .B(AB[1]), .C(n1331[0]), 
         .D(n1331[1]), .Z(n20883)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(B (D)))) */ ;   // c:/s_links/sources/quad_decoder.v(106[36:38])
    defparam i15940_4_lut_4_lut_4_lut.init = 16'h6620;
    LUT4 mux_859_i25_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[24]), 
         .D(quad_count_adj_529[24]), .Z(\spi_data_out_r_39__N_1547[24] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i15_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[14]), 
         .D(quad_count_adj_531[14]), .Z(\spi_data_out_r_39__N_2249[14] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i22_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[21]), 
         .D(quad_count_adj_533[21]), .Z(\spi_data_out_r_39__N_2015[21] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i21_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[20]), 
         .D(quad_count_adj_533[20]), .Z(\spi_data_out_r_39__N_2015[20] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i14_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[13]), 
         .D(quad_count_adj_531[13]), .Z(\spi_data_out_r_39__N_2249[13] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i20_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[19]), 
         .D(quad_count_adj_533[19]), .Z(\spi_data_out_r_39__N_2015[19] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i19_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[18]), 
         .D(quad_count_adj_533[18]), .Z(\spi_data_out_r_39__N_2015[18] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i18_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[17]), 
         .D(quad_count_adj_533[17]), .Z(\spi_data_out_r_39__N_2015[17] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i13_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[12]), 
         .D(quad_count_adj_531[12]), .Z(\spi_data_out_r_39__N_2249[12] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i17_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[16]), 
         .D(quad_count_adj_533[16]), .Z(\spi_data_out_r_39__N_2015[16] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i16_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[15]), 
         .D(quad_count_adj_533[15]), .Z(\spi_data_out_r_39__N_2015[15] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i15_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[14]), 
         .D(quad_count_adj_533[14]), .Z(\spi_data_out_r_39__N_2015[14] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i14_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[13]), 
         .D(quad_count_adj_533[13]), .Z(\spi_data_out_r_39__N_2015[13] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i12_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[11]), 
         .D(quad_count_adj_531[11]), .Z(\spi_data_out_r_39__N_2249[11] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i11_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[10]), 
         .D(quad_count_adj_531[10]), .Z(\spi_data_out_r_39__N_2249[10] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i10_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[9]), 
         .D(quad_count_adj_531[9]), .Z(\spi_data_out_r_39__N_2249[9] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i10_3_lut_4_lut.init = 16'hf1e0;
    FD1S3IX i41_407 (.D(spi_data_out_r_39__N_1162), .CK(clk), .CD(n29239), 
            .Q(spi_data_out_r_39__N_974)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam i41_407.GSR = "DISABLED";
    LUT4 mux_862_i9_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[8]), 
         .D(quad_count_adj_531[8]), .Z(\spi_data_out_r_39__N_2249[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i9_3_lut_4_lut.init = 16'hf1e0;
    FD1S3IX quad_set_complete_451 (.D(quad_set_valid), .CK(clk_1MHz), .CD(n29239), 
            .Q(quad_set_complete)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_set_complete_451.GSR = "DISABLED";
    LUT4 mux_861_i13_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[12]), 
         .D(quad_count_adj_533[12]), .Z(\spi_data_out_r_39__N_2015[12] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i12_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[11]), 
         .D(quad_count_adj_533[11]), .Z(\spi_data_out_r_39__N_2015[11] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i8_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[7]), 
         .D(quad_count_adj_531[7]), .Z(\spi_data_out_r_39__N_2249[7] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i7_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[6]), 
         .D(quad_count_adj_531[6]), .Z(\spi_data_out_r_39__N_2249[6] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i6_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[5]), 
         .D(quad_count_adj_531[5]), .Z(\spi_data_out_r_39__N_2249[5] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i5_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[4]), 
         .D(quad_count_adj_531[4]), .Z(\spi_data_out_r_39__N_2249[4] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i24_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[23]), 
         .D(quad_count_adj_529[23]), .Z(\spi_data_out_r_39__N_1547[23] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i11_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[10]), 
         .D(quad_count_adj_533[10]), .Z(\spi_data_out_r_39__N_2015[10] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i10_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[9]), 
         .D(quad_count_adj_533[9]), .Z(\spi_data_out_r_39__N_2015[9] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i4_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[3]), 
         .D(quad_count_adj_531[3]), .Z(\spi_data_out_r_39__N_2249[3] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i9_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[8]), 
         .D(quad_count_adj_533[8]), .Z(\spi_data_out_r_39__N_2015[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i8_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[7]), 
         .D(quad_count_adj_533[7]), .Z(\spi_data_out_r_39__N_2015[7] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i7_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[6]), 
         .D(quad_count_adj_533[6]), .Z(\spi_data_out_r_39__N_2015[6] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i6_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[5]), 
         .D(quad_count_adj_533[5]), .Z(\spi_data_out_r_39__N_2015[5] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i23_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[22]), 
         .D(quad_count_adj_529[22]), .Z(\spi_data_out_r_39__N_1547[22] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i3_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[2]), 
         .D(quad_count_adj_531[2]), .Z(\spi_data_out_r_39__N_2249[2] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i22_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[21]), 
         .D(quad_count_adj_529[21]), .Z(\spi_data_out_r_39__N_1547[21] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i5_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[4]), 
         .D(quad_count_adj_533[4]), .Z(\spi_data_out_r_39__N_2015[4] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i4_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[3]), 
         .D(quad_count_adj_533[3]), .Z(\spi_data_out_r_39__N_2015[3] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i21_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[20]), 
         .D(quad_count_adj_529[20]), .Z(\spi_data_out_r_39__N_1547[20] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_862_i2_3_lut_4_lut (.A(n29098), .B(n13511), .C(quad_buffer_adj_530[1]), 
         .D(quad_count_adj_531[1]), .Z(\spi_data_out_r_39__N_2249[1] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_862_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i3_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[2]), 
         .D(quad_count_adj_533[2]), .Z(\spi_data_out_r_39__N_2015[2] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i2_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[1]), 
         .D(quad_count_adj_533[1]), .Z(\spi_data_out_r_39__N_2015[1] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i1_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[0]), 
         .D(quad_count_adj_535[0]), .Z(\spi_data_out_r_39__N_1781[0] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i20_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[19]), 
         .D(quad_count_adj_529[19]), .Z(\spi_data_out_r_39__N_1547[19] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i32_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[31]), 
         .D(quad_count_adj_535[31]), .Z(\spi_data_out_r_39__N_1781[31] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i31_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[30]), 
         .D(quad_count_adj_535[30]), .Z(\spi_data_out_r_39__N_1781[30] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i30_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[29]), 
         .D(quad_count_adj_535[29]), .Z(\spi_data_out_r_39__N_1781[29] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i29_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[28]), 
         .D(quad_count_adj_535[28]), .Z(\spi_data_out_r_39__N_1781[28] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i28_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[27]), 
         .D(quad_count_adj_535[27]), .Z(\spi_data_out_r_39__N_1781[27] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_531 (.A(n1331[1]), .B(n1331[2]), .Z(n29259)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_531.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_944 (.A(n1331[1]), .B(n1331[2]), .C(AB[0]), 
         .Z(n4)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_944.init = 16'he0e0;
    LUT4 i117_2_lut_3_lut_4_lut (.A(quad_homing[1]), .B(quad_homing[0]), 
         .C(n29260), .D(pin_io_out_4), .Z(n108)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam i117_2_lut_3_lut_4_lut.init = 16'hfbff;
    LUT4 i1_2_lut_3_lut_4_lut (.A(quad_homing[1]), .B(quad_homing[0]), .C(n29260), 
         .D(pin_io_out_4), .Z(n79)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0400;
    LUT4 mux_860_i27_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[26]), 
         .D(quad_count_adj_535[26]), .Z(\spi_data_out_r_39__N_1781[26] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i19_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[18]), 
         .D(quad_count_adj_529[18]), .Z(\spi_data_out_r_39__N_1547[18] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i18_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[17]), 
         .D(quad_count_adj_529[17]), .Z(\spi_data_out_r_39__N_1547[17] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i26_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[25]), 
         .D(quad_count_adj_535[25]), .Z(\spi_data_out_r_39__N_1781[25] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i25_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[24]), 
         .D(quad_count_adj_535[24]), .Z(\spi_data_out_r_39__N_1781[24] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i24_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[23]), 
         .D(quad_count_adj_535[23]), .Z(\spi_data_out_r_39__N_1781[23] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i42_2_lut_rep_533 (.A(AB[0]), .B(AB[1]), .Z(n29261)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(106[36:38])
    defparam i42_2_lut_rep_533.init = 16'h6666;
    LUT4 mux_859_i17_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[16]), 
         .D(quad_count_adj_529[16]), .Z(\spi_data_out_r_39__N_1547[16] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i32_4_lut_4_lut (.A(AB[0]), .B(AB[1]), .C(n4), .D(n1331[3]), 
         .Z(n9539)) /* synthesis lut_function=(A (B (C+(D)))+!A !(B ((D)+!C)+!B !(D))) */ ;   // c:/s_links/sources/quad_decoder.v(106[36:38])
    defparam i32_4_lut_4_lut.init = 16'h99c0;
    LUT4 mux_860_i23_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[22]), 
         .D(quad_count_adj_535[22]), .Z(\spi_data_out_r_39__N_1781[22] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i22_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[21]), 
         .D(quad_count_adj_535[21]), .Z(\spi_data_out_r_39__N_1781[21] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i21_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[20]), 
         .D(quad_count_adj_535[20]), .Z(\spi_data_out_r_39__N_1781[20] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i20_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[19]), 
         .D(quad_count_adj_535[19]), .Z(\spi_data_out_r_39__N_1781[19] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i19_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[18]), 
         .D(quad_count_adj_535[18]), .Z(\spi_data_out_r_39__N_1781[18] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i16_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[15]), 
         .D(quad_count_adj_529[15]), .Z(\spi_data_out_r_39__N_1547[15] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i15_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[14]), 
         .D(quad_count_adj_529[14]), .Z(\spi_data_out_r_39__N_1547[14] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i18_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[17]), 
         .D(quad_count_adj_535[17]), .Z(\spi_data_out_r_39__N_1781[17] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i17_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[16]), 
         .D(quad_count_adj_535[16]), .Z(\spi_data_out_r_39__N_1781[16] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n100_bdd_4_lut (.A(n29259), .B(n1331[0]), .C(AB[0]), .D(AB[1]), 
         .Z(n29034)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D)))) */ ;
    defparam n100_bdd_4_lut.init = 16'hc00e;
    LUT4 mux_860_i16_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[15]), 
         .D(quad_count_adj_535[15]), .Z(\spi_data_out_r_39__N_1781[15] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i15_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[14]), 
         .D(quad_count_adj_535[14]), .Z(\spi_data_out_r_39__N_1781[14] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i14_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[13]), 
         .D(quad_count_adj_535[13]), .Z(\spi_data_out_r_39__N_1781[13] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i13_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[12]), 
         .D(quad_count_adj_535[12]), .Z(\spi_data_out_r_39__N_1781[12] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i12_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[11]), 
         .D(quad_count_adj_535[11]), .Z(\spi_data_out_r_39__N_1781[11] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i12_3_lut_4_lut.init = 16'hf1e0;
    FD1S3IX state_FSM_i3 (.D(n9539), .CK(clk_1MHz), .CD(n29239), .Q(n1331[3]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i3.GSR = "DISABLED";
    FD1S3IX state_FSM_i2 (.D(n29322), .CK(clk_1MHz), .CD(n29239), .Q(n1331[2]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i2.GSR = "DISABLED";
    FD1S3IX state_FSM_i1 (.D(n9547), .CK(clk_1MHz), .CD(n29239), .Q(n1331[1]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i1.GSR = "DISABLED";
    LUT4 mux_859_i14_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[13]), 
         .D(quad_count_adj_529[13]), .Z(\spi_data_out_r_39__N_1547[13] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i11_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[10]), 
         .D(quad_count_adj_535[10]), .Z(\spi_data_out_r_39__N_1781[10] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i10_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[9]), 
         .D(quad_count_adj_535[9]), .Z(\spi_data_out_r_39__N_1781[9] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i9_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[8]), 
         .D(quad_count_adj_535[8]), .Z(\spi_data_out_r_39__N_1781[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i8_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[7]), 
         .D(quad_count_adj_535[7]), .Z(\spi_data_out_r_39__N_1781[7] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i7_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[6]), 
         .D(quad_count_adj_535[6]), .Z(\spi_data_out_r_39__N_1781[6] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i6_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[5]), 
         .D(quad_count_adj_535[5]), .Z(\spi_data_out_r_39__N_1781[5] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_3_lut_4_lut (.A(n27256), .B(n29078), .C(n27338), .D(n29213), 
         .Z(clk_enable_199)) /* synthesis lut_function=(A (B (C+!(D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h8088;
    LUT4 mux_860_i5_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[4]), 
         .D(quad_count_adj_535[4]), .Z(\spi_data_out_r_39__N_1781[4] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i4_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[3]), 
         .D(quad_count_adj_535[3]), .Z(\spi_data_out_r_39__N_1781[3] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i3_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[2]), 
         .D(quad_count_adj_535[2]), .Z(\spi_data_out_r_39__N_1781[2] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_860_i2_3_lut_4_lut (.A(n13413), .B(n29098), .C(quad_buffer_adj_534[1]), 
         .D(quad_count_adj_535[1]), .Z(\spi_data_out_r_39__N_1781[1] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_860_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_863_i1_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[0]), 
         .D(quad_count[0]), .Z(\spi_data_out_r_39__N_2483[0] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i32_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[31]), 
         .D(quad_count[31]), .Z(\spi_data_out_r_39__N_2483[31] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i32_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i39_4_lut (.A(AB[0]), .B(AB[1]), .C(n1331[2]), .D(n1331[1]), 
         .Z(n51)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C+(D)))+!A (B+!(C)))) */ ;
    defparam i39_4_lut.init = 16'h1812;
    LUT4 mux_863_i31_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[30]), 
         .D(quad_count[30]), .Z(\spi_data_out_r_39__N_2483[30] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i31_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i30_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[29]), 
         .D(quad_count[29]), .Z(\spi_data_out_r_39__N_2483[29] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i30_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i29_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[28]), 
         .D(quad_count[28]), .Z(\spi_data_out_r_39__N_2483[28] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i29_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_859_i1_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[0]), 
         .D(quad_count_adj_529[0]), .Z(\spi_data_out_r_39__N_1547[0] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_863_i28_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[27]), 
         .D(quad_count[27]), .Z(\spi_data_out_r_39__N_2483[27] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i28_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i27_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[26]), 
         .D(quad_count[26]), .Z(\spi_data_out_r_39__N_2483[26] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i27_3_lut_4_lut.init = 16'hf4b0;
    CCU2D add_2145_33 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[30]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[31]), 
          .D1(GND_net), .CIN(n25070), .S0(n6496[30]), .S1(n6496[31]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_33.INIT0 = 16'h7878;
    defparam add_2145_33.INIT1 = 16'h7878;
    defparam add_2145_33.INJECT1_0 = "NO";
    defparam add_2145_33.INJECT1_1 = "NO";
    LUT4 mux_863_i26_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[25]), 
         .D(quad_count[25]), .Z(\spi_data_out_r_39__N_2483[25] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i26_3_lut_4_lut.init = 16'hf4b0;
    CCU2D add_2145_31 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[28]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[29]), 
          .D1(GND_net), .CIN(n25069), .COUT(n25070), .S0(n6496[28]), 
          .S1(n6496[29]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_31.INIT0 = 16'h7878;
    defparam add_2145_31.INIT1 = 16'h7878;
    defparam add_2145_31.INJECT1_0 = "NO";
    defparam add_2145_31.INJECT1_1 = "NO";
    CCU2D add_2145_29 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[26]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[27]), 
          .D1(GND_net), .CIN(n25068), .COUT(n25069), .S0(n6496[26]), 
          .S1(n6496[27]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_29.INIT0 = 16'h7878;
    defparam add_2145_29.INIT1 = 16'h7878;
    defparam add_2145_29.INJECT1_0 = "NO";
    defparam add_2145_29.INJECT1_1 = "NO";
    CCU2D add_2145_27 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[24]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[25]), 
          .D1(GND_net), .CIN(n25067), .COUT(n25068), .S0(n6496[24]), 
          .S1(n6496[25]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_27.INIT0 = 16'h7878;
    defparam add_2145_27.INIT1 = 16'h7878;
    defparam add_2145_27.INJECT1_0 = "NO";
    defparam add_2145_27.INJECT1_1 = "NO";
    CCU2D add_2145_25 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[22]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[23]), 
          .D1(GND_net), .CIN(n25066), .COUT(n25067), .S0(n6496[22]), 
          .S1(n6496[23]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_25.INIT0 = 16'h7878;
    defparam add_2145_25.INIT1 = 16'h7878;
    defparam add_2145_25.INJECT1_0 = "NO";
    defparam add_2145_25.INJECT1_1 = "NO";
    CCU2D add_2145_23 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[20]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[21]), 
          .D1(GND_net), .CIN(n25065), .COUT(n25066), .S0(n6496[20]), 
          .S1(n6496[21]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_23.INIT0 = 16'h7878;
    defparam add_2145_23.INIT1 = 16'h7878;
    defparam add_2145_23.INJECT1_0 = "NO";
    defparam add_2145_23.INJECT1_1 = "NO";
    CCU2D add_2145_21 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[18]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[19]), 
          .D1(GND_net), .CIN(n25064), .COUT(n25065), .S0(n6496[18]), 
          .S1(n6496[19]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_21.INIT0 = 16'h7878;
    defparam add_2145_21.INIT1 = 16'h7878;
    defparam add_2145_21.INJECT1_0 = "NO";
    defparam add_2145_21.INJECT1_1 = "NO";
    CCU2D add_2145_19 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[16]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[17]), 
          .D1(GND_net), .CIN(n25063), .COUT(n25064), .S0(n6496[16]), 
          .S1(n6496[17]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_19.INIT0 = 16'h7878;
    defparam add_2145_19.INIT1 = 16'h7878;
    defparam add_2145_19.INJECT1_0 = "NO";
    defparam add_2145_19.INJECT1_1 = "NO";
    CCU2D add_2145_17 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[14]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[15]), 
          .D1(GND_net), .CIN(n25062), .COUT(n25063), .S0(n6496[14]), 
          .S1(n6496[15]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_17.INIT0 = 16'h7878;
    defparam add_2145_17.INIT1 = 16'h7878;
    defparam add_2145_17.INJECT1_0 = "NO";
    defparam add_2145_17.INJECT1_1 = "NO";
    CCU2D add_2145_15 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[12]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[13]), 
          .D1(GND_net), .CIN(n25061), .COUT(n25062), .S0(n6496[12]), 
          .S1(n6496[13]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_15.INIT0 = 16'h7878;
    defparam add_2145_15.INIT1 = 16'h7878;
    defparam add_2145_15.INJECT1_0 = "NO";
    defparam add_2145_15.INJECT1_1 = "NO";
    LUT4 mux_863_i25_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[24]), 
         .D(quad_count[24]), .Z(\spi_data_out_r_39__N_2483[24] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i25_3_lut_4_lut.init = 16'hf4b0;
    CCU2D add_2145_13 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[10]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[11]), 
          .D1(GND_net), .CIN(n25060), .COUT(n25061), .S0(n6496[10]), 
          .S1(n6496[11]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_13.INIT0 = 16'h7878;
    defparam add_2145_13.INIT1 = 16'h7878;
    defparam add_2145_13.INJECT1_0 = "NO";
    defparam add_2145_13.INJECT1_1 = "NO";
    LUT4 mux_863_i24_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[23]), 
         .D(quad_count[23]), .Z(\spi_data_out_r_39__N_2483[23] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i24_3_lut_4_lut.init = 16'hf4b0;
    CCU2D add_2145_11 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[8]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[9]), 
          .D1(GND_net), .CIN(n25059), .COUT(n25060), .S0(n6496[8]), 
          .S1(n6496[9]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_11.INIT0 = 16'h7878;
    defparam add_2145_11.INIT1 = 16'h7878;
    defparam add_2145_11.INJECT1_0 = "NO";
    defparam add_2145_11.INJECT1_1 = "NO";
    CCU2D add_2145_9 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[6]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[7]), 
          .D1(GND_net), .CIN(n25058), .COUT(n25059), .S0(n6496[6]), 
          .S1(n6496[7]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_9.INIT0 = 16'h7878;
    defparam add_2145_9.INIT1 = 16'h7878;
    defparam add_2145_9.INJECT1_0 = "NO";
    defparam add_2145_9.INJECT1_1 = "NO";
    LUT4 mux_863_i23_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[22]), 
         .D(quad_count[22]), .Z(\spi_data_out_r_39__N_2483[22] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i23_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i22_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[21]), 
         .D(quad_count[21]), .Z(\spi_data_out_r_39__N_2483[21] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i22_3_lut_4_lut.init = 16'hf4b0;
    CCU2D add_2145_7 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[4]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[5]), 
          .D1(GND_net), .CIN(n25057), .COUT(n25058), .S0(n6496[4]), 
          .S1(n6496[5]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_7.INIT0 = 16'h7878;
    defparam add_2145_7.INIT1 = 16'h7878;
    defparam add_2145_7.INJECT1_0 = "NO";
    defparam add_2145_7.INJECT1_1 = "NO";
    CCU2D add_2145_5 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[2]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[3]), 
          .D1(GND_net), .CIN(n25056), .COUT(n25057), .S0(n6496[2]), 
          .S1(n6496[3]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_5.INIT0 = 16'h7878;
    defparam add_2145_5.INIT1 = 16'h7878;
    defparam add_2145_5.INJECT1_0 = "NO";
    defparam add_2145_5.INJECT1_1 = "NO";
    CCU2D add_2145_3 (.A0(resetn_c), .B0(n41), .C0(quad_count_adj_7594[0]), 
          .D0(GND_net), .A1(resetn_c), .B1(n41), .C1(quad_count_adj_7594[1]), 
          .D1(GND_net), .CIN(n25055), .COUT(n25056), .S0(n6496[0]), 
          .S1(n6496[1]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_3.INIT0 = 16'h8787;
    defparam add_2145_3.INIT1 = 16'h7878;
    defparam add_2145_3.INJECT1_0 = "NO";
    defparam add_2145_3.INJECT1_1 = "NO";
    CCU2D add_2145_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(resetn_c), .B1(n41), .C1(GND_net), .D1(GND_net), .COUT(n25055));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2145_1.INIT0 = 16'hF000;
    defparam add_2145_1.INIT1 = 16'h7777;
    defparam add_2145_1.INJECT1_0 = "NO";
    defparam add_2145_1.INJECT1_1 = "NO";
    LUT4 mux_863_i21_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[20]), 
         .D(quad_count[20]), .Z(\spi_data_out_r_39__N_2483[20] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i21_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i20_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[19]), 
         .D(quad_count[19]), .Z(\spi_data_out_r_39__N_2483[19] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i20_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i19_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[18]), 
         .D(quad_count[18]), .Z(\spi_data_out_r_39__N_2483[18] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i19_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i18_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[17]), 
         .D(quad_count[17]), .Z(\spi_data_out_r_39__N_2483[17] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i18_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_859_i13_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[12]), 
         .D(quad_count_adj_529[12]), .Z(\spi_data_out_r_39__N_1547[12] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_863_i17_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[16]), 
         .D(quad_count[16]), .Z(\spi_data_out_r_39__N_2483[16] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i17_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_859_i32_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[31]), 
         .D(quad_count_adj_529[31]), .Z(\spi_data_out_r_39__N_1547[31] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_863_i16_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[15]), 
         .D(quad_count[15]), .Z(\spi_data_out_r_39__N_2483[15] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i16_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_859_i31_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[30]), 
         .D(quad_count_adj_529[30]), .Z(\spi_data_out_r_39__N_1547[30] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_863_i15_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[14]), 
         .D(quad_count[14]), .Z(\spi_data_out_r_39__N_2483[14] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i15_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_859_i12_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[11]), 
         .D(quad_count_adj_529[11]), .Z(\spi_data_out_r_39__N_1547[11] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i11_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[10]), 
         .D(quad_count_adj_529[10]), .Z(\spi_data_out_r_39__N_1547[10] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_863_i14_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[13]), 
         .D(quad_count[13]), .Z(\spi_data_out_r_39__N_2483[13] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i14_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_859_i10_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[9]), 
         .D(quad_count_adj_529[9]), .Z(\spi_data_out_r_39__N_1547[9] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i37_4_lut_else_3_lut (.A(n1331[2]), .B(AB[0]), .C(AB[1]), .D(n1331[0]), 
         .Z(n29320)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C (D))))) */ ;
    defparam i37_4_lut_else_3_lut.init = 16'h3828;
    LUT4 mux_863_i13_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[12]), 
         .D(quad_count[12]), .Z(\spi_data_out_r_39__N_2483[12] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i13_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i12_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[11]), 
         .D(quad_count[11]), .Z(\spi_data_out_r_39__N_2483[11] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i12_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_863_i11_3_lut_4_lut (.A(n29099), .B(n25293), .C(quad_buffer[10]), 
         .D(quad_count[10]), .Z(\spi_data_out_r_39__N_2483[10] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_863_i11_3_lut_4_lut.init = 16'hf4b0;
    FD1S3AX quad_buffer_i31 (.D(quad_count_adj_7594[31]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i31.GSR = "DISABLED";
    FD1S3AX quad_buffer_i30 (.D(quad_count_adj_7594[30]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i30.GSR = "DISABLED";
    FD1S3AX quad_buffer_i29 (.D(quad_count_adj_7594[29]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i29.GSR = "DISABLED";
    FD1S3AX quad_buffer_i28 (.D(quad_count_adj_7594[28]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i28.GSR = "DISABLED";
    FD1S3AX quad_buffer_i27 (.D(quad_count_adj_7594[27]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i27.GSR = "DISABLED";
    FD1S3AX quad_buffer_i26 (.D(quad_count_adj_7594[26]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i26.GSR = "DISABLED";
    FD1S3AX quad_buffer_i25 (.D(quad_count_adj_7594[25]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i25.GSR = "DISABLED";
    FD1S3AX quad_buffer_i24 (.D(quad_count_adj_7594[24]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i24.GSR = "DISABLED";
    FD1S3AX quad_buffer_i23 (.D(quad_count_adj_7594[23]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i23.GSR = "DISABLED";
    FD1S3AX quad_buffer_i22 (.D(quad_count_adj_7594[22]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i22.GSR = "DISABLED";
    FD1S3AX quad_buffer_i21 (.D(quad_count_adj_7594[21]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i21.GSR = "DISABLED";
    FD1S3AX quad_buffer_i20 (.D(quad_count_adj_7594[20]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i20.GSR = "DISABLED";
    FD1S3AX quad_buffer_i19 (.D(quad_count_adj_7594[19]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i19.GSR = "DISABLED";
    FD1S3AX quad_buffer_i18 (.D(quad_count_adj_7594[18]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i18.GSR = "DISABLED";
    FD1S3AX quad_buffer_i17 (.D(quad_count_adj_7594[17]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i17.GSR = "DISABLED";
    FD1S3AX quad_buffer_i16 (.D(quad_count_adj_7594[16]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i16.GSR = "DISABLED";
    FD1S3AX quad_buffer_i15 (.D(quad_count_adj_7594[15]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i15.GSR = "DISABLED";
    FD1S3AX quad_buffer_i14 (.D(quad_count_adj_7594[14]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i14.GSR = "DISABLED";
    FD1S3AX quad_buffer_i13 (.D(quad_count_adj_7594[13]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i13.GSR = "DISABLED";
    FD1S3AX quad_buffer_i12 (.D(quad_count_adj_7594[12]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i12.GSR = "DISABLED";
    FD1S3AX quad_buffer_i11 (.D(quad_count_adj_7594[11]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i11.GSR = "DISABLED";
    FD1S3AX quad_buffer_i10 (.D(quad_count_adj_7594[10]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i10.GSR = "DISABLED";
    FD1S3AX quad_buffer_i9 (.D(quad_count_adj_7594[9]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i9.GSR = "DISABLED";
    FD1S3AX quad_buffer_i8 (.D(quad_count_adj_7594[8]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i8.GSR = "DISABLED";
    FD1S3AX quad_buffer_i7 (.D(quad_count_adj_7594[7]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i7.GSR = "DISABLED";
    FD1S3AX quad_buffer_i6 (.D(quad_count_adj_7594[6]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i6.GSR = "DISABLED";
    FD1S3AX quad_buffer_i5 (.D(quad_count_adj_7594[5]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i5.GSR = "DISABLED";
    FD1S3AX quad_buffer_i4 (.D(quad_count_adj_7594[4]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i4.GSR = "DISABLED";
    FD1S3AX quad_buffer_i3 (.D(quad_count_adj_7594[3]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i3.GSR = "DISABLED";
    FD1S3AX quad_buffer_i2 (.D(quad_count_adj_7594[2]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i2.GSR = "DISABLED";
    FD1S3AX quad_buffer_i1 (.D(quad_count_adj_7594[1]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer_adj_7595[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i1.GSR = "DISABLED";
    FD1S3AX AB_i1 (.D(sync[1]), .CK(clk_1MHz), .Q(AB[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam AB_i1.GSR = "DISABLED";
    LUT4 mux_859_i9_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[8]), 
         .D(quad_count_adj_529[8]), .Z(\spi_data_out_r_39__N_1547[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2_3_lut (.A(\spi_addr[1] ), .B(\spi_addr[2] ), .C(n29761), .Z(n25293)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_3_lut.init = 16'h8080;
    FD1S3AX sync_i1 (.D(\quad_a[0] ), .CK(clk_1MHz), .Q(sync[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam sync_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(spi_data_out_r_39__N_1079[31]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i31 (.D(spi_data_out_r_39__N_1079[30]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i30 (.D(spi_data_out_r_39__N_1079[29]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    LUT4 mux_859_i8_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[7]), 
         .D(quad_count_adj_529[7]), .Z(\spi_data_out_r_39__N_1547[7] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i8_3_lut_4_lut.init = 16'hf1e0;
    FD1S3AX spi_data_out_r_i29 (.D(spi_data_out_r_39__N_1079[28]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i28 (.D(spi_data_out_r_39__N_1079[27]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i27 (.D(spi_data_out_r_39__N_1079[26]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i26 (.D(spi_data_out_r_39__N_1079[25]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i25 (.D(spi_data_out_r_39__N_1079[24]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i24 (.D(spi_data_out_r_39__N_1079[23]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i23 (.D(spi_data_out_r_39__N_1079[22]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i22 (.D(spi_data_out_r_39__N_1079[21]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i21 (.D(spi_data_out_r_39__N_1079[20]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i20 (.D(spi_data_out_r_39__N_1079[19]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i19 (.D(spi_data_out_r_39__N_1079[18]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i18 (.D(spi_data_out_r_39__N_1079[17]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i17 (.D(spi_data_out_r_39__N_1079[16]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i16 (.D(spi_data_out_r_39__N_1079[15]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(spi_data_out_r_39__N_1079[14]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(spi_data_out_r_39__N_1079[13]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(spi_data_out_r_39__N_1079[12]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(spi_data_out_r_39__N_1079[11]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(spi_data_out_r_39__N_1079[10]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(spi_data_out_r_39__N_1079[9]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(spi_data_out_r_39__N_1079[8]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(spi_data_out_r_39__N_1079[7]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(spi_data_out_r_39__N_1079[6]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(spi_data_out_r_39__N_1079[5]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(spi_data_out_r_39__N_1079[4]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(spi_data_out_r_39__N_1079[3]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(spi_data_out_r_39__N_1079[2]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(spi_data_out_r_39__N_1079[1]), .CK(clk), 
            .Q(\spi_data_out_r_39__N_934[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    LUT4 mux_859_i7_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[6]), 
         .D(quad_count_adj_529[6]), .Z(\spi_data_out_r_39__N_1547[6] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i7_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX quad_count_i0_i31 (.D(n10353), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i31.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i30 (.D(n10355), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i30.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i29 (.D(n10357), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i29.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i28 (.D(n10359), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i28.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i27 (.D(n10361), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i27.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i26 (.D(n10363), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i26.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i25 (.D(n10365), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i25.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i24 (.D(n10367), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i24.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i23 (.D(n10369), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i23.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i22 (.D(n10371), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i22.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i21 (.D(n10373), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i21.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i20 (.D(n10375), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i20.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i19 (.D(n10377), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i19.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i18 (.D(n10379), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i18.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i17 (.D(n10381), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i17.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i16 (.D(n10383), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i16.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i15 (.D(n10385), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i15.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i14 (.D(n10387), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i14.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i13 (.D(n10389), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i13.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i12 (.D(n10391), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i12.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i11 (.D(n10393), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i11.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i10 (.D(n10395), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i10.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i9 (.D(n10397), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i9.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i8 (.D(n10399), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i8.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i7 (.D(n10401), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i7.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i6 (.D(n10403), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i6.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i5 (.D(n10405), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i5.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i4 (.D(n10407), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i4.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i3 (.D(n10409), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i3.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i2 (.D(n10411), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i1 (.D(n10413), .SP(clk_1MHz_enable_340), .CK(clk_1MHz), 
            .Q(quad_count_adj_7594[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i1.GSR = "DISABLED";
    LUT4 mux_859_i6_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[5]), 
         .D(quad_count_adj_529[5]), .Z(\spi_data_out_r_39__N_1547[5] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i5_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[4]), 
         .D(quad_count_adj_529[4]), .Z(\spi_data_out_r_39__N_1547[4] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i4_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[3]), 
         .D(quad_count_adj_529[3]), .Z(\spi_data_out_r_39__N_1547[3] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i3_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[2]), 
         .D(quad_count_adj_529[2]), .Z(\spi_data_out_r_39__N_1547[2] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_859_i2_3_lut_4_lut (.A(n13413), .B(n29099), .C(quad_buffer_adj_528[1]), 
         .D(quad_count_adj_529[1]), .Z(\spi_data_out_r_39__N_1547[1] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_859_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i1_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[0]), 
         .D(quad_count_adj_537[0]), .Z(\spi_data_out_r_39__N_1313[0] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i32_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[31]), 
         .D(quad_count_adj_537[31]), .Z(\spi_data_out_r_39__N_1313[31] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i22901_3_lut_4_lut (.A(\spi_cmd[2] ), .B(n29117), .C(\spi_addr[2] ), 
         .D(n29310), .Z(clear_intrpt_N_3065)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam i22901_3_lut_4_lut.init = 16'h0010;
    LUT4 mux_858_i31_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[30]), 
         .D(quad_count_adj_537[30]), .Z(\spi_data_out_r_39__N_1313[30] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i30_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[29]), 
         .D(quad_count_adj_537[29]), .Z(\spi_data_out_r_39__N_1313[29] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i29_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[28]), 
         .D(quad_count_adj_537[28]), .Z(\spi_data_out_r_39__N_1313[28] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i28_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[27]), 
         .D(quad_count_adj_537[27]), .Z(\spi_data_out_r_39__N_1313[27] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i28_3_lut_4_lut.init = 16'hf1e0;
    FD1P3IX quad_set__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i1.GSR = "DISABLED";
    FD1P3IX quad_set__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i2.GSR = "DISABLED";
    FD1P3IX quad_set__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i3.GSR = "DISABLED";
    FD1P3IX quad_set__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i4.GSR = "DISABLED";
    FD1P3IX quad_set__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i5.GSR = "DISABLED";
    FD1P3IX quad_set__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i6.GSR = "DISABLED";
    FD1P3IX quad_set__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i7.GSR = "DISABLED";
    FD1P3IX quad_set__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i8.GSR = "DISABLED";
    FD1P3IX quad_set__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i9.GSR = "DISABLED";
    FD1P3IX quad_set__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i10.GSR = "DISABLED";
    FD1P3IX quad_set__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i11.GSR = "DISABLED";
    FD1P3IX quad_set__i12 (.D(\spi_data_r[12] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i12.GSR = "DISABLED";
    FD1P3IX quad_set__i13 (.D(\spi_data_r[13] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i13.GSR = "DISABLED";
    FD1P3IX quad_set__i14 (.D(\spi_data_r[14] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i14.GSR = "DISABLED";
    FD1P3IX quad_set__i15 (.D(\spi_data_r[15] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i15.GSR = "DISABLED";
    FD1P3IX quad_set__i16 (.D(\spi_data_r[16] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i16.GSR = "DISABLED";
    FD1P3IX quad_set__i17 (.D(\spi_data_r[17] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i17.GSR = "DISABLED";
    FD1P3IX quad_set__i18 (.D(\spi_data_r[18] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i18.GSR = "DISABLED";
    FD1P3IX quad_set__i19 (.D(\spi_data_r[19] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i19.GSR = "DISABLED";
    FD1P3IX quad_set__i20 (.D(\spi_data_r[20] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i20.GSR = "DISABLED";
    FD1P3IX quad_set__i21 (.D(\spi_data_r[21] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i21.GSR = "DISABLED";
    FD1P3IX quad_set__i22 (.D(\spi_data_r[22] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i22.GSR = "DISABLED";
    FD1P3IX quad_set__i23 (.D(\spi_data_r[23] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i23.GSR = "DISABLED";
    FD1P3IX quad_set__i24 (.D(\spi_data_r[24] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i24.GSR = "DISABLED";
    FD1P3IX quad_set__i25 (.D(\spi_data_r[25] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i25.GSR = "DISABLED";
    FD1P3IX quad_set__i26 (.D(\spi_data_r[26] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i26.GSR = "DISABLED";
    FD1P3IX quad_set__i27 (.D(\spi_data_r[27] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i27.GSR = "DISABLED";
    FD1P3IX quad_set__i28 (.D(\spi_data_r[28] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i28.GSR = "DISABLED";
    FD1P3IX quad_set__i29 (.D(\spi_data_r[29] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i29.GSR = "DISABLED";
    FD1P3IX quad_set__i30 (.D(\spi_data_r[30] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i30.GSR = "DISABLED";
    FD1P3IX quad_set__i31 (.D(\spi_data_r[31] ), .SP(clk_enable_433), .CD(n29239), 
            .CK(clk), .Q(quad_set[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i31.GSR = "DISABLED";
    FD1P3IX quad_homing__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_436), .CD(n29239), 
            .CK(clk), .Q(quad_homing[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam quad_homing__i1.GSR = "DISABLED";
    FD1P3IX quad_set_valid_404 (.D(n29085), .SP(clk_enable_501), .CD(n29239), 
            .CK(clk), .Q(quad_set_valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set_valid_404.GSR = "DISABLED";
    LUT4 mux_858_i27_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[26]), 
         .D(quad_count_adj_537[26]), .Z(\spi_data_out_r_39__N_1313[26] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i26_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[25]), 
         .D(quad_count_adj_537[25]), .Z(\spi_data_out_r_39__N_1313[25] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i25_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[24]), 
         .D(quad_count_adj_537[24]), .Z(\spi_data_out_r_39__N_1313[24] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5560_4_lut (.A(n6496[31]), .B(quad_set[31]), .C(n3), .D(n26), 
         .Z(n10353)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5560_4_lut.init = 16'hc0ca;
    LUT4 i5562_4_lut (.A(n6496[30]), .B(quad_set[30]), .C(n3), .D(n26), 
         .Z(n10355)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5562_4_lut.init = 16'hc0ca;
    LUT4 i5564_4_lut (.A(n6496[29]), .B(quad_set[29]), .C(n3), .D(n26), 
         .Z(n10357)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5564_4_lut.init = 16'hc0ca;
    LUT4 i5566_4_lut (.A(n6496[28]), .B(quad_set[28]), .C(n3), .D(n26), 
         .Z(n10359)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5566_4_lut.init = 16'hc0ca;
    LUT4 i5568_4_lut (.A(n6496[27]), .B(quad_set[27]), .C(n3), .D(n26), 
         .Z(n10361)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5568_4_lut.init = 16'hc0ca;
    LUT4 i5570_4_lut (.A(n6496[26]), .B(quad_set[26]), .C(n3), .D(n26), 
         .Z(n10363)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5570_4_lut.init = 16'hc0ca;
    LUT4 i5572_4_lut (.A(n6496[25]), .B(quad_set[25]), .C(n3), .D(n26), 
         .Z(n10365)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5572_4_lut.init = 16'hc0ca;
    LUT4 i5574_4_lut (.A(n6496[24]), .B(quad_set[24]), .C(n3), .D(n26), 
         .Z(n10367)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5574_4_lut.init = 16'hc0ca;
    LUT4 i5576_4_lut (.A(n6496[23]), .B(quad_set[23]), .C(n3), .D(n26), 
         .Z(n10369)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5576_4_lut.init = 16'hc0ca;
    LUT4 i5578_4_lut (.A(n6496[22]), .B(quad_set[22]), .C(n3), .D(n26), 
         .Z(n10371)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5578_4_lut.init = 16'hc0ca;
    LUT4 mux_858_i24_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[23]), 
         .D(quad_count_adj_537[23]), .Z(\spi_data_out_r_39__N_1313[23] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5580_4_lut (.A(n6496[21]), .B(quad_set[21]), .C(n3), .D(n26), 
         .Z(n10373)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5580_4_lut.init = 16'hc0ca;
    LUT4 mux_858_i23_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[22]), 
         .D(quad_count_adj_537[22]), .Z(\spi_data_out_r_39__N_1313[22] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i22_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[21]), 
         .D(quad_count_adj_537[21]), .Z(\spi_data_out_r_39__N_1313[21] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i21_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[20]), 
         .D(quad_count_adj_537[20]), .Z(\spi_data_out_r_39__N_1313[20] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i20_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[19]), 
         .D(quad_count_adj_537[19]), .Z(\spi_data_out_r_39__N_1313[19] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i19_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[18]), 
         .D(quad_count_adj_537[18]), .Z(\spi_data_out_r_39__N_1313[18] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5582_4_lut (.A(n6496[20]), .B(quad_set[20]), .C(n3), .D(n26), 
         .Z(n10375)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5582_4_lut.init = 16'hc0ca;
    LUT4 i5584_4_lut (.A(n6496[19]), .B(quad_set[19]), .C(n3), .D(n26), 
         .Z(n10377)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5584_4_lut.init = 16'hc0ca;
    LUT4 i5586_4_lut (.A(n6496[18]), .B(quad_set[18]), .C(n3), .D(n26), 
         .Z(n10379)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5586_4_lut.init = 16'hc0ca;
    LUT4 i5588_4_lut (.A(n6496[17]), .B(quad_set[17]), .C(n3), .D(n26), 
         .Z(n10381)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5588_4_lut.init = 16'hc0ca;
    LUT4 i5590_4_lut (.A(n6496[16]), .B(quad_set[16]), .C(n3), .D(n26), 
         .Z(n10383)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5590_4_lut.init = 16'hc0ca;
    LUT4 i5592_4_lut (.A(n6496[15]), .B(quad_set[15]), .C(n3), .D(n26), 
         .Z(n10385)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5592_4_lut.init = 16'hc0ca;
    LUT4 i5594_4_lut (.A(n6496[14]), .B(quad_set[14]), .C(n3), .D(n26), 
         .Z(n10387)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5594_4_lut.init = 16'hc0ca;
    LUT4 i5596_4_lut (.A(n6496[13]), .B(quad_set[13]), .C(n3), .D(n26), 
         .Z(n10389)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5596_4_lut.init = 16'hc0ca;
    LUT4 i5598_4_lut (.A(n6496[12]), .B(quad_set[12]), .C(n3), .D(n26), 
         .Z(n10391)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5598_4_lut.init = 16'hc0ca;
    LUT4 i5600_4_lut (.A(n6496[11]), .B(quad_set[11]), .C(n3), .D(n26), 
         .Z(n10393)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5600_4_lut.init = 16'hc0ca;
    LUT4 i5602_4_lut (.A(n6496[10]), .B(quad_set[10]), .C(n3), .D(n26), 
         .Z(n10395)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5602_4_lut.init = 16'hc0ca;
    LUT4 i5604_4_lut (.A(n6496[9]), .B(quad_set[9]), .C(n3), .D(n26), 
         .Z(n10397)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5604_4_lut.init = 16'hc0ca;
    LUT4 i5606_4_lut (.A(n6496[8]), .B(quad_set[8]), .C(n3), .D(n26), 
         .Z(n10399)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5606_4_lut.init = 16'hc0ca;
    LUT4 i5608_4_lut (.A(n6496[7]), .B(quad_set[7]), .C(n3), .D(n26), 
         .Z(n10401)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5608_4_lut.init = 16'hc0ca;
    LUT4 i5610_4_lut (.A(n6496[6]), .B(quad_set[6]), .C(n3), .D(n26), 
         .Z(n10403)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5610_4_lut.init = 16'hc0ca;
    LUT4 i5612_4_lut (.A(n6496[5]), .B(quad_set[5]), .C(n3), .D(n26), 
         .Z(n10405)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5612_4_lut.init = 16'hc0ca;
    LUT4 mux_858_i18_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[17]), 
         .D(quad_count_adj_537[17]), .Z(\spi_data_out_r_39__N_1313[17] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i5614_4_lut (.A(n6496[4]), .B(quad_set[4]), .C(n3), .D(n26), 
         .Z(n10407)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5614_4_lut.init = 16'hc0ca;
    LUT4 i5616_4_lut (.A(n6496[3]), .B(quad_set[3]), .C(n3), .D(n26), 
         .Z(n10409)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5616_4_lut.init = 16'hc0ca;
    LUT4 i5618_4_lut (.A(n6496[2]), .B(quad_set[2]), .C(n3), .D(n26), 
         .Z(n10411)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5618_4_lut.init = 16'hc0ca;
    LUT4 i5620_4_lut (.A(n6496[1]), .B(quad_set[1]), .C(n3), .D(n26), 
         .Z(n10413)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5620_4_lut.init = 16'hc0ca;
    LUT4 i15876_4_lut (.A(n1331[2]), .B(n29261), .C(n1331[1]), .D(n1331[3]), 
         .Z(n20819)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;
    defparam i15876_4_lut.init = 16'hcc36;
    LUT4 mux_858_i17_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[16]), 
         .D(quad_count_adj_537[16]), .Z(\spi_data_out_r_39__N_1313[16] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i4670_4_lut (.A(n6496[0]), .B(quad_set[0]), .C(n3), .D(n26), 
         .Z(n9438)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i4670_4_lut.init = 16'hc0ca;
    LUT4 mux_858_i16_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[15]), 
         .D(quad_count_adj_537[15]), .Z(\spi_data_out_r_39__N_1313[15] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i15_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[14]), 
         .D(quad_count_adj_537[14]), .Z(\spi_data_out_r_39__N_1313[14] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i49_4_lut (.A(n1331[2]), .B(n1331[3]), .C(n1331[1]), .D(n29261), 
         .Z(n31)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (D)+!B !(C (D)+!C !(D))))) */ ;
    defparam i49_4_lut.init = 16'h32cd;
    LUT4 mux_858_i14_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[13]), 
         .D(quad_count_adj_537[13]), .Z(\spi_data_out_r_39__N_1313[13] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i13_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[12]), 
         .D(quad_count_adj_537[12]), .Z(\spi_data_out_r_39__N_1313[12] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i12_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[11]), 
         .D(quad_count_adj_537[11]), .Z(\spi_data_out_r_39__N_1313[11] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i11_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[10]), 
         .D(quad_count_adj_537[10]), .Z(\spi_data_out_r_39__N_1313[10] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i10_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[9]), 
         .D(quad_count_adj_537[9]), .Z(\spi_data_out_r_39__N_1313[9] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i9_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[8]), 
         .D(quad_count_adj_537[8]), .Z(\spi_data_out_r_39__N_1313[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i8_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[7]), 
         .D(quad_count_adj_537[7]), .Z(\spi_data_out_r_39__N_1313[7] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i7_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[6]), 
         .D(quad_count_adj_537[6]), .Z(\spi_data_out_r_39__N_1313[6] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i6_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[5]), 
         .D(quad_count_adj_537[5]), .Z(\spi_data_out_r_39__N_1313[5] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i5_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[4]), 
         .D(quad_count_adj_537[4]), .Z(\spi_data_out_r_39__N_1313[4] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i4_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[3]), 
         .D(quad_count_adj_537[3]), .Z(\spi_data_out_r_39__N_1313[3] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i3_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[2]), 
         .D(quad_count_adj_537[2]), .Z(\spi_data_out_r_39__N_1313[2] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_858_i2_3_lut_4_lut (.A(n29098), .B(n13506), .C(quad_buffer_adj_536[1]), 
         .D(quad_count_adj_537[1]), .Z(\spi_data_out_r_39__N_1313[1] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_858_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i1_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[0]), 
         .D(quad_count_adj_7594[0]), .Z(spi_data_out_r_39__N_1079[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i32_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[31]), 
         .D(quad_count_adj_7594[31]), .Z(spi_data_out_r_39__N_1079[31])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i31_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[30]), 
         .D(quad_count_adj_7594[30]), .Z(spi_data_out_r_39__N_1079[30])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i30_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[29]), 
         .D(quad_count_adj_7594[29]), .Z(spi_data_out_r_39__N_1079[29])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i29_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[28]), 
         .D(quad_count_adj_7594[28]), .Z(spi_data_out_r_39__N_1079[28])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i29_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i28_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[27]), 
         .D(quad_count_adj_7594[27]), .Z(spi_data_out_r_39__N_1079[27])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i28_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i27_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[26]), 
         .D(quad_count_adj_7594[26]), .Z(spi_data_out_r_39__N_1079[26])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i27_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i26_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[25]), 
         .D(quad_count_adj_7594[25]), .Z(spi_data_out_r_39__N_1079[25])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i26_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i25_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[24]), 
         .D(quad_count_adj_7594[24]), .Z(spi_data_out_r_39__N_1079[24])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i25_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i24_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[23]), 
         .D(quad_count_adj_7594[23]), .Z(spi_data_out_r_39__N_1079[23])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i24_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i23_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[22]), 
         .D(quad_count_adj_7594[22]), .Z(spi_data_out_r_39__N_1079[22])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i23_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i22_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[21]), 
         .D(quad_count_adj_7594[21]), .Z(spi_data_out_r_39__N_1079[21])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i22_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i21_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[20]), 
         .D(quad_count_adj_7594[20]), .Z(spi_data_out_r_39__N_1079[20])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i21_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i20_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[19]), 
         .D(quad_count_adj_7594[19]), .Z(spi_data_out_r_39__N_1079[19])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i20_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i19_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[18]), 
         .D(quad_count_adj_7594[18]), .Z(spi_data_out_r_39__N_1079[18])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i19_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i18_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[17]), 
         .D(quad_count_adj_7594[17]), .Z(spi_data_out_r_39__N_1079[17])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i18_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i17_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[16]), 
         .D(quad_count_adj_7594[16]), .Z(spi_data_out_r_39__N_1079[16])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i17_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i16_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[15]), 
         .D(quad_count_adj_7594[15]), .Z(spi_data_out_r_39__N_1079[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i15_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[14]), 
         .D(quad_count_adj_7594[14]), .Z(spi_data_out_r_39__N_1079[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i14_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[13]), 
         .D(quad_count_adj_7594[13]), .Z(spi_data_out_r_39__N_1079[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i14_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i13_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[12]), 
         .D(quad_count_adj_7594[12]), .Z(spi_data_out_r_39__N_1079[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i12_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[11]), 
         .D(quad_count_adj_7594[11]), .Z(spi_data_out_r_39__N_1079[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i12_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i23156 (.BLUT(n29320), .ALUT(n29321), .C0(n1331[3]), .Z(n29322));
    LUT4 mux_857_i11_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[10]), 
         .D(quad_count_adj_7594[10]), .Z(spi_data_out_r_39__N_1079[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i10_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[9]), 
         .D(quad_count_adj_7594[9]), .Z(spi_data_out_r_39__N_1079[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i9_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[8]), 
         .D(quad_count_adj_7594[8]), .Z(spi_data_out_r_39__N_1079[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i8_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[7]), 
         .D(quad_count_adj_7594[7]), .Z(spi_data_out_r_39__N_1079[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i7_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[6]), 
         .D(quad_count_adj_7594[6]), .Z(spi_data_out_r_39__N_1079[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i6_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[5]), 
         .D(quad_count_adj_7594[5]), .Z(spi_data_out_r_39__N_1079[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i5_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[4]), 
         .D(quad_count_adj_7594[4]), .Z(spi_data_out_r_39__N_1079[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i4_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[3]), 
         .D(quad_count_adj_7594[3]), .Z(spi_data_out_r_39__N_1079[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_4_lut (.A(n20883), .B(AB[1]), .C(AB[0]), .D(n1331[3]), .Z(n9547)) /* synthesis lut_function=(A+!(B+!(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hbaaa;
    LUT4 mux_857_i3_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[2]), 
         .D(quad_count_adj_7594[2]), .Z(spi_data_out_r_39__N_1079[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i1_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[0]), 
         .D(quad_count_adj_533[0]), .Z(\spi_data_out_r_39__N_2015[0] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_857_i2_3_lut_4_lut (.A(n29099), .B(n13506), .C(quad_buffer_adj_7595[1]), 
         .D(quad_count_adj_7594[1]), .Z(spi_data_out_r_39__N_1079[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_857_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i32_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[31]), 
         .D(quad_count_adj_533[31]), .Z(\spi_data_out_r_39__N_2015[31] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i32_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i31_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[30]), 
         .D(quad_count_adj_533[30]), .Z(\spi_data_out_r_39__N_2015[30] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i31_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_861_i30_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[29]), 
         .D(quad_count_adj_533[29]), .Z(\spi_data_out_r_39__N_2015[29] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i30_3_lut_4_lut.init = 16'hf1e0;
    LUT4 AB_0__bdd_4_lut_23253 (.A(AB[0]), .B(n29259), .C(n1331[3]), .D(AB[1]), 
         .Z(n29326)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(B (C (D)+!C !(D))+!B (D))) */ ;
    defparam AB_0__bdd_4_lut_23253.init = 16'ha659;
    LUT4 mux_861_i29_3_lut_4_lut (.A(n29099), .B(n13511), .C(quad_buffer_adj_532[28]), 
         .D(quad_count_adj_533[28]), .Z(\spi_data_out_r_39__N_2015[28] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(78[11:41])
    defparam mux_861_i29_3_lut_4_lut.init = 16'hf1e0;
    
endmodule
//
// Verilog Description of module \quad_decoder(DEV_ID=2) 
//

module \quad_decoder(DEV_ID=2)  (quad_count, clk_1MHz, \spi_data_out_r_39__N_1402[0] , 
            clk, \spi_data_out_r_39__N_1547[0] , \quad_b[2] , quad_buffer, 
            \mode[2]_derived_32 , clk_enable_269, n29239, \spi_data_r[0] , 
            n26948, quad_homing, clk_enable_435, n29762, spi_data_out_r_39__N_1442, 
            quad_set_complete, n29099, \spi_addr[0] , n26933, n13506, 
            spi_data_out_r_39__N_1162, n13413, resetn_c, n13511, spi_data_out_r_39__N_2098, 
            n25293, spi_data_out_r_39__N_2566, pin_io_out_24, n29233, 
            \spi_data_r[31] , \spi_data_r[30] , \spi_data_r[29] , \spi_data_r[28] , 
            \spi_data_r[27] , \spi_data_r[26] , \spi_data_r[25] , \spi_data_r[24] , 
            \spi_data_r[23] , \spi_data_r[22] , \spi_data_r[21] , \spi_data_r[20] , 
            \spi_data_r[19] , \spi_data_r[18] , \spi_data_r[17] , \spi_data_r[16] , 
            \spi_data_r[15] , \spi_data_r[14] , \spi_data_r[13] , \spi_data_r[12] , 
            \spi_data_r[11] , \spi_data_r[10] , \spi_data_r[9] , \spi_data_r[8] , 
            \spi_data_r[7] , \spi_data_r[6] , \spi_data_r[5] , \spi_data_r[4] , 
            \spi_data_r[3] , \spi_data_r[2] , \spi_data_r[1] , \quad_a[2] , 
            \spi_data_out_r_39__N_1402[31] , \spi_data_out_r_39__N_1547[31] , 
            \spi_data_out_r_39__N_1402[30] , \spi_data_out_r_39__N_1547[30] , 
            \spi_data_out_r_39__N_1402[29] , \spi_data_out_r_39__N_1547[29] , 
            \spi_data_out_r_39__N_1402[28] , \spi_data_out_r_39__N_1547[28] , 
            \spi_data_out_r_39__N_1402[27] , \spi_data_out_r_39__N_1547[27] , 
            \spi_data_out_r_39__N_1402[26] , \spi_data_out_r_39__N_1547[26] , 
            \spi_data_out_r_39__N_1402[25] , \spi_data_out_r_39__N_1547[25] , 
            \spi_data_out_r_39__N_1402[24] , \spi_data_out_r_39__N_1547[24] , 
            \spi_data_out_r_39__N_1402[23] , \spi_data_out_r_39__N_1547[23] , 
            \spi_data_out_r_39__N_1402[22] , \spi_data_out_r_39__N_1547[22] , 
            \spi_data_out_r_39__N_1402[21] , \spi_data_out_r_39__N_1547[21] , 
            \spi_data_out_r_39__N_1402[20] , \spi_data_out_r_39__N_1547[20] , 
            \spi_data_out_r_39__N_1402[19] , \spi_data_out_r_39__N_1547[19] , 
            \spi_data_out_r_39__N_1402[18] , \spi_data_out_r_39__N_1547[18] , 
            \spi_data_out_r_39__N_1402[17] , \spi_data_out_r_39__N_1547[17] , 
            \spi_data_out_r_39__N_1402[16] , \spi_data_out_r_39__N_1547[16] , 
            \spi_data_out_r_39__N_1402[15] , \spi_data_out_r_39__N_1547[15] , 
            \spi_data_out_r_39__N_1402[14] , \spi_data_out_r_39__N_1547[14] , 
            \spi_data_out_r_39__N_1402[13] , \spi_data_out_r_39__N_1547[13] , 
            \spi_data_out_r_39__N_1402[12] , \spi_data_out_r_39__N_1547[12] , 
            \spi_data_out_r_39__N_1402[11] , \spi_data_out_r_39__N_1547[11] , 
            \spi_data_out_r_39__N_1402[10] , \spi_data_out_r_39__N_1547[10] , 
            \spi_data_out_r_39__N_1402[9] , \spi_data_out_r_39__N_1547[9] , 
            \spi_data_out_r_39__N_1402[8] , \spi_data_out_r_39__N_1547[8] , 
            \spi_data_out_r_39__N_1402[7] , \spi_data_out_r_39__N_1547[7] , 
            \spi_data_out_r_39__N_1402[6] , \spi_data_out_r_39__N_1547[6] , 
            \spi_data_out_r_39__N_1402[5] , \spi_data_out_r_39__N_1547[5] , 
            \spi_data_out_r_39__N_1402[4] , \spi_data_out_r_39__N_1547[4] , 
            \spi_data_out_r_39__N_1402[3] , \spi_data_out_r_39__N_1547[3] , 
            \spi_data_out_r_39__N_1402[2] , \spi_data_out_r_39__N_1547[2] , 
            \spi_data_out_r_39__N_1402[1] , \spi_data_out_r_39__N_1547[1] , 
            n27301, clk_enable_503, n29122, GND_net, n29326, n108, 
            quad_set_valid, n3, mem_rdata_update_N_729, n9633, n12714, 
            n13, n29336, n95, quad_set_valid_adj_207, n5647) /* synthesis syn_module_defined=1 */ ;
    output [31:0]quad_count;
    input clk_1MHz;
    output \spi_data_out_r_39__N_1402[0] ;
    input clk;
    input \spi_data_out_r_39__N_1547[0] ;
    input \quad_b[2] ;
    output [31:0]quad_buffer;
    input \mode[2]_derived_32 ;
    input clk_enable_269;
    input n29239;
    input \spi_data_r[0] ;
    output n26948;
    output [1:0]quad_homing;
    input clk_enable_435;
    input n29762;
    output spi_data_out_r_39__N_1442;
    output quad_set_complete;
    input n29099;
    input \spi_addr[0] ;
    input n26933;
    input n13506;
    output spi_data_out_r_39__N_1162;
    input n13413;
    input resetn_c;
    input n13511;
    output spi_data_out_r_39__N_2098;
    input n25293;
    output spi_data_out_r_39__N_2566;
    input pin_io_out_24;
    input n29233;
    input \spi_data_r[31] ;
    input \spi_data_r[30] ;
    input \spi_data_r[29] ;
    input \spi_data_r[28] ;
    input \spi_data_r[27] ;
    input \spi_data_r[26] ;
    input \spi_data_r[25] ;
    input \spi_data_r[24] ;
    input \spi_data_r[23] ;
    input \spi_data_r[22] ;
    input \spi_data_r[21] ;
    input \spi_data_r[20] ;
    input \spi_data_r[19] ;
    input \spi_data_r[18] ;
    input \spi_data_r[17] ;
    input \spi_data_r[16] ;
    input \spi_data_r[15] ;
    input \spi_data_r[14] ;
    input \spi_data_r[13] ;
    input \spi_data_r[12] ;
    input \spi_data_r[11] ;
    input \spi_data_r[10] ;
    input \spi_data_r[9] ;
    input \spi_data_r[8] ;
    input \spi_data_r[7] ;
    input \spi_data_r[6] ;
    input \spi_data_r[5] ;
    input \spi_data_r[4] ;
    input \spi_data_r[3] ;
    input \spi_data_r[2] ;
    input \spi_data_r[1] ;
    input \quad_a[2] ;
    output \spi_data_out_r_39__N_1402[31] ;
    input \spi_data_out_r_39__N_1547[31] ;
    output \spi_data_out_r_39__N_1402[30] ;
    input \spi_data_out_r_39__N_1547[30] ;
    output \spi_data_out_r_39__N_1402[29] ;
    input \spi_data_out_r_39__N_1547[29] ;
    output \spi_data_out_r_39__N_1402[28] ;
    input \spi_data_out_r_39__N_1547[28] ;
    output \spi_data_out_r_39__N_1402[27] ;
    input \spi_data_out_r_39__N_1547[27] ;
    output \spi_data_out_r_39__N_1402[26] ;
    input \spi_data_out_r_39__N_1547[26] ;
    output \spi_data_out_r_39__N_1402[25] ;
    input \spi_data_out_r_39__N_1547[25] ;
    output \spi_data_out_r_39__N_1402[24] ;
    input \spi_data_out_r_39__N_1547[24] ;
    output \spi_data_out_r_39__N_1402[23] ;
    input \spi_data_out_r_39__N_1547[23] ;
    output \spi_data_out_r_39__N_1402[22] ;
    input \spi_data_out_r_39__N_1547[22] ;
    output \spi_data_out_r_39__N_1402[21] ;
    input \spi_data_out_r_39__N_1547[21] ;
    output \spi_data_out_r_39__N_1402[20] ;
    input \spi_data_out_r_39__N_1547[20] ;
    output \spi_data_out_r_39__N_1402[19] ;
    input \spi_data_out_r_39__N_1547[19] ;
    output \spi_data_out_r_39__N_1402[18] ;
    input \spi_data_out_r_39__N_1547[18] ;
    output \spi_data_out_r_39__N_1402[17] ;
    input \spi_data_out_r_39__N_1547[17] ;
    output \spi_data_out_r_39__N_1402[16] ;
    input \spi_data_out_r_39__N_1547[16] ;
    output \spi_data_out_r_39__N_1402[15] ;
    input \spi_data_out_r_39__N_1547[15] ;
    output \spi_data_out_r_39__N_1402[14] ;
    input \spi_data_out_r_39__N_1547[14] ;
    output \spi_data_out_r_39__N_1402[13] ;
    input \spi_data_out_r_39__N_1547[13] ;
    output \spi_data_out_r_39__N_1402[12] ;
    input \spi_data_out_r_39__N_1547[12] ;
    output \spi_data_out_r_39__N_1402[11] ;
    input \spi_data_out_r_39__N_1547[11] ;
    output \spi_data_out_r_39__N_1402[10] ;
    input \spi_data_out_r_39__N_1547[10] ;
    output \spi_data_out_r_39__N_1402[9] ;
    input \spi_data_out_r_39__N_1547[9] ;
    output \spi_data_out_r_39__N_1402[8] ;
    input \spi_data_out_r_39__N_1547[8] ;
    output \spi_data_out_r_39__N_1402[7] ;
    input \spi_data_out_r_39__N_1547[7] ;
    output \spi_data_out_r_39__N_1402[6] ;
    input \spi_data_out_r_39__N_1547[6] ;
    output \spi_data_out_r_39__N_1402[5] ;
    input \spi_data_out_r_39__N_1547[5] ;
    output \spi_data_out_r_39__N_1402[4] ;
    input \spi_data_out_r_39__N_1547[4] ;
    output \spi_data_out_r_39__N_1402[3] ;
    input \spi_data_out_r_39__N_1547[3] ;
    output \spi_data_out_r_39__N_1402[2] ;
    input \spi_data_out_r_39__N_1547[2] ;
    output \spi_data_out_r_39__N_1402[1] ;
    input \spi_data_out_r_39__N_1547[1] ;
    input n27301;
    input clk_enable_503;
    input n29122;
    input GND_net;
    input n29326;
    input n108;
    input quad_set_valid;
    output n3;
    input mem_rdata_update_N_729;
    output n9633;
    input n12714;
    output n13;
    input n29336;
    input n95;
    input quad_set_valid_adj_207;
    output n5647;
    
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire [1:0]sync /* synthesis ASYNC_REG="TRUE" */ ;   // c:/s_links/sources/quad_decoder.v(106[30:34])
    wire [1:0]AB /* synthesis ASYNC_REG="TRUE" */ ;   // c:/s_links/sources/quad_decoder.v(106[36:38])
    wire \mode[2]_derived_32  /* synthesis is_clock=1, SET_AS_NETWORK=\stepper_ins[2].u_stepper/mode[2]_derived_32 */ ;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    
    wire clk_1MHz_enable_278, n14;
    wire [31:0]quad_set;   // c:/s_links/sources/quad_decoder.v(40[31:39])
    wire [3:0]n1711;
    
    wire n28870, n11568, n11606, n29234, n6, n26795, n9470, n59, 
        n26751, spi_data_out_r_39__N_1630, quad_set_valid_c, n28607, 
        n29053, n36, n14_adj_7176, n14_adj_7177, n14_adj_7178, n14_adj_7179, 
        n14_adj_7180, n14_adj_7181, n14_adj_7182, n14_adj_7183, n14_adj_7184, 
        n14_adj_7185, n14_adj_7186, n14_adj_7187, n14_adj_7188, n14_adj_7189, 
        n14_adj_7190, n14_adj_7191, n14_adj_7192, n14_adj_7193, n14_adj_7194, 
        n14_adj_7195, n14_adj_7196, n14_adj_7197, n14_adj_7198, n14_adj_7199, 
        n14_adj_7200, n14_adj_7201, n14_adj_7202, n14_adj_7203, n14_adj_7204, 
        n14_adj_7205, n14_adj_7206;
    wire [31:0]n6301;
    
    wire n3_c, n25150, n25149, n25148, n25147, n25146, n25145, 
        n25144, n25143, n25142, n25141, n25140, n25139, n25138, 
        n25137, n25136, n25135, n12820;
    
    FD1P3AX quad_count_i0_i0 (.D(n14), .SP(clk_1MHz_enable_278), .CK(clk_1MHz), 
            .Q(quad_count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_1547[0] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX sync_i0 (.D(\quad_b[2] ), .CK(clk_1MHz), .Q(sync[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam sync_i0.GSR = "DISABLED";
    FD1S3AX AB_i0 (.D(sync[0]), .CK(clk_1MHz), .Q(AB[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam AB_i0.GSR = "DISABLED";
    FD1S3AX quad_buffer_i0 (.D(quad_count[0]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i0.GSR = "DISABLED";
    FD1P3IX quad_set__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i0.GSR = "DISABLED";
    FD1S3JX state_FSM_i0 (.D(n28870), .CK(clk_1MHz), .PD(n29239), .Q(n1711[0]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i0.GSR = "DISABLED";
    LUT4 i4672_3_lut_4_lut (.A(AB[0]), .B(AB[1]), .C(n1711[3]), .D(n11568), 
         .Z(n11606)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // c:/s_links/sources/quad_decoder.v(162[19:30])
    defparam i4672_3_lut_4_lut.init = 16'hbfb0;
    LUT4 i15_2_lut_rep_506 (.A(AB[1]), .B(AB[0]), .Z(n29234)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(155[16] 158[10])
    defparam i15_2_lut_rep_506.init = 16'h6666;
    LUT4 i1_3_lut_4_lut (.A(AB[1]), .B(AB[0]), .C(n1711[2]), .D(n1711[3]), 
         .Z(n26948)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(D))) */ ;   // c:/s_links/sources/quad_decoder.v(155[16] 158[10])
    defparam i1_3_lut_4_lut.init = 16'h9960;
    LUT4 i1_4_lut_4_lut (.A(AB[1]), .B(AB[0]), .C(n1711[1]), .D(n6), 
         .Z(n26795)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C+(D))))) */ ;   // c:/s_links/sources/quad_decoder.v(155[16] 158[10])
    defparam i1_4_lut_4_lut.init = 16'h6460;
    FD1P3IX quad_homing__i0 (.D(n29762), .SP(clk_enable_435), .CD(n29239), 
            .CK(clk), .Q(quad_homing[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam quad_homing__i0.GSR = "DISABLED";
    LUT4 i4697_4_lut_4_lut (.A(n1711[2]), .B(AB[0]), .C(AB[1]), .D(n6), 
         .Z(n9470)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C (D))))) */ ;   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam i4697_4_lut_4_lut.init = 16'h3828;
    LUT4 i1_4_lut_4_lut_adj_906 (.A(n1711[3]), .B(AB[0]), .C(AB[1]), .D(n59), 
         .Z(n26751)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i1_4_lut_4_lut_adj_906.init = 16'h96c3;
    FD1S3IX i41_407 (.D(spi_data_out_r_39__N_1630), .CK(clk), .CD(n29239), 
            .Q(spi_data_out_r_39__N_1442)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam i41_407.GSR = "DISABLED";
    FD1S3IX quad_set_complete_451 (.D(quad_set_valid_c), .CK(clk_1MHz), 
            .CD(n29239), .Q(quad_set_complete)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_set_complete_451.GSR = "DISABLED";
    LUT4 n59_bdd_4_lut_23102 (.A(n59), .B(n1711[3]), .C(AB[1]), .D(AB[0]), 
         .Z(n28607)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C (D)))+!A (B (C (D)+!C !(D)))) */ ;
    defparam n59_bdd_4_lut_23102.init = 16'he00c;
    LUT4 i22586_2_lut_2_lut_4_lut (.A(n29099), .B(\spi_addr[0] ), .C(n26933), 
         .D(n13506), .Z(spi_data_out_r_39__N_1162)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (D))) */ ;
    defparam i22586_2_lut_2_lut_4_lut.init = 16'h0057;
    LUT4 i22595_2_lut_2_lut_4_lut (.A(n29099), .B(\spi_addr[0] ), .C(n26933), 
         .D(n13413), .Z(spi_data_out_r_39__N_1630)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (D))) */ ;
    defparam i22595_2_lut_2_lut_4_lut.init = 16'h0057;
    LUT4 n1712_bdd_4_lut (.A(n1711[3]), .B(n29234), .C(n1711[2]), .D(resetn_c), 
         .Z(n29053)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C (D))))) */ ;
    defparam n1712_bdd_4_lut.init = 16'h6200;
    LUT4 i22604_2_lut_2_lut_4_lut (.A(n29099), .B(\spi_addr[0] ), .C(n26933), 
         .D(n13511), .Z(spi_data_out_r_39__N_2098)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (D))) */ ;
    defparam i22604_2_lut_2_lut_4_lut.init = 16'h0057;
    LUT4 i22612_2_lut_2_lut_4_lut (.A(n29099), .B(\spi_addr[0] ), .C(n26933), 
         .D(n25293), .Z(spi_data_out_r_39__N_2566)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(D))) */ ;
    defparam i22612_2_lut_2_lut_4_lut.init = 16'h5700;
    FD1S3IX state_FSM_i3 (.D(n28607), .CK(clk_1MHz), .CD(n29239), .Q(n1711[3]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i3.GSR = "DISABLED";
    FD1S3IX state_FSM_i2 (.D(n9470), .CK(clk_1MHz), .CD(n29239), .Q(n1711[2]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i2.GSR = "DISABLED";
    FD1S3IX state_FSM_i1 (.D(n26795), .CK(clk_1MHz), .CD(n29239), .Q(n1711[1]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i1.GSR = "DISABLED";
    LUT4 i3_3_lut_4_lut (.A(pin_io_out_24), .B(n29233), .C(quad_homing[0]), 
         .D(quad_homing[1]), .Z(n36)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i3_3_lut_4_lut.init = 16'hffdf;
    FD1P3IX quad_set__i31 (.D(\spi_data_r[31] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i31.GSR = "DISABLED";
    FD1P3IX quad_set__i30 (.D(\spi_data_r[30] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i30.GSR = "DISABLED";
    FD1P3IX quad_set__i29 (.D(\spi_data_r[29] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i29.GSR = "DISABLED";
    FD1P3IX quad_set__i28 (.D(\spi_data_r[28] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i28.GSR = "DISABLED";
    FD1P3IX quad_set__i27 (.D(\spi_data_r[27] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i27.GSR = "DISABLED";
    FD1P3IX quad_set__i26 (.D(\spi_data_r[26] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i26.GSR = "DISABLED";
    FD1P3IX quad_set__i25 (.D(\spi_data_r[25] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i25.GSR = "DISABLED";
    FD1P3IX quad_set__i24 (.D(\spi_data_r[24] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i24.GSR = "DISABLED";
    FD1P3IX quad_set__i23 (.D(\spi_data_r[23] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i23.GSR = "DISABLED";
    FD1P3IX quad_set__i22 (.D(\spi_data_r[22] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i22.GSR = "DISABLED";
    FD1P3IX quad_set__i21 (.D(\spi_data_r[21] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i21.GSR = "DISABLED";
    FD1P3IX quad_set__i20 (.D(\spi_data_r[20] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i20.GSR = "DISABLED";
    FD1P3IX quad_set__i19 (.D(\spi_data_r[19] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i19.GSR = "DISABLED";
    FD1P3IX quad_set__i18 (.D(\spi_data_r[18] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i18.GSR = "DISABLED";
    FD1P3IX quad_set__i17 (.D(\spi_data_r[17] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i17.GSR = "DISABLED";
    FD1P3IX quad_set__i16 (.D(\spi_data_r[16] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i16.GSR = "DISABLED";
    FD1P3IX quad_set__i15 (.D(\spi_data_r[15] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i15.GSR = "DISABLED";
    FD1P3IX quad_set__i14 (.D(\spi_data_r[14] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i14.GSR = "DISABLED";
    FD1P3IX quad_set__i13 (.D(\spi_data_r[13] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i13.GSR = "DISABLED";
    FD1P3IX quad_set__i12 (.D(\spi_data_r[12] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i12.GSR = "DISABLED";
    FD1P3IX quad_set__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i11.GSR = "DISABLED";
    FD1P3IX quad_set__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i10.GSR = "DISABLED";
    FD1P3IX quad_set__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i9.GSR = "DISABLED";
    FD1P3IX quad_set__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i8.GSR = "DISABLED";
    FD1P3IX quad_set__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i7.GSR = "DISABLED";
    FD1P3IX quad_set__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i6.GSR = "DISABLED";
    FD1P3IX quad_set__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i5.GSR = "DISABLED";
    FD1P3IX quad_set__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i4.GSR = "DISABLED";
    FD1P3IX quad_set__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i3.GSR = "DISABLED";
    FD1P3IX quad_set__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i2.GSR = "DISABLED";
    FD1P3IX quad_set__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_269), .CD(n29239), 
            .CK(clk), .Q(quad_set[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i1.GSR = "DISABLED";
    LUT4 i4671_4_lut (.A(AB[0]), .B(AB[1]), .C(n1711[2]), .D(n1711[1]), 
         .Z(n11568)) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A (B+!(C))) */ ;
    defparam i4671_4_lut.init = 16'he7ed;
    FD1S3AX quad_buffer_i31 (.D(quad_count[31]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i31.GSR = "DISABLED";
    FD1S3AX quad_buffer_i30 (.D(quad_count[30]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i30.GSR = "DISABLED";
    FD1S3AX quad_buffer_i29 (.D(quad_count[29]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i29.GSR = "DISABLED";
    FD1S3AX quad_buffer_i28 (.D(quad_count[28]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i28.GSR = "DISABLED";
    FD1S3AX quad_buffer_i27 (.D(quad_count[27]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i27.GSR = "DISABLED";
    FD1S3AX quad_buffer_i26 (.D(quad_count[26]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i26.GSR = "DISABLED";
    FD1S3AX quad_buffer_i25 (.D(quad_count[25]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i25.GSR = "DISABLED";
    FD1S3AX quad_buffer_i24 (.D(quad_count[24]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i24.GSR = "DISABLED";
    FD1S3AX quad_buffer_i23 (.D(quad_count[23]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i23.GSR = "DISABLED";
    FD1S3AX quad_buffer_i22 (.D(quad_count[22]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i22.GSR = "DISABLED";
    FD1S3AX quad_buffer_i21 (.D(quad_count[21]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i21.GSR = "DISABLED";
    FD1S3AX quad_buffer_i20 (.D(quad_count[20]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i20.GSR = "DISABLED";
    FD1S3AX quad_buffer_i19 (.D(quad_count[19]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i19.GSR = "DISABLED";
    FD1S3AX quad_buffer_i18 (.D(quad_count[18]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i18.GSR = "DISABLED";
    FD1S3AX quad_buffer_i17 (.D(quad_count[17]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i17.GSR = "DISABLED";
    FD1S3AX quad_buffer_i16 (.D(quad_count[16]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i16.GSR = "DISABLED";
    FD1S3AX quad_buffer_i15 (.D(quad_count[15]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i15.GSR = "DISABLED";
    FD1S3AX quad_buffer_i14 (.D(quad_count[14]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i14.GSR = "DISABLED";
    FD1S3AX quad_buffer_i13 (.D(quad_count[13]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i13.GSR = "DISABLED";
    FD1S3AX quad_buffer_i12 (.D(quad_count[12]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i12.GSR = "DISABLED";
    FD1S3AX quad_buffer_i11 (.D(quad_count[11]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i11.GSR = "DISABLED";
    FD1S3AX quad_buffer_i10 (.D(quad_count[10]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i10.GSR = "DISABLED";
    FD1S3AX quad_buffer_i9 (.D(quad_count[9]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i9.GSR = "DISABLED";
    FD1S3AX quad_buffer_i8 (.D(quad_count[8]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i8.GSR = "DISABLED";
    FD1S3AX quad_buffer_i7 (.D(quad_count[7]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i7.GSR = "DISABLED";
    FD1S3AX quad_buffer_i6 (.D(quad_count[6]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i6.GSR = "DISABLED";
    FD1S3AX quad_buffer_i5 (.D(quad_count[5]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i5.GSR = "DISABLED";
    FD1S3AX quad_buffer_i4 (.D(quad_count[4]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i4.GSR = "DISABLED";
    FD1S3AX quad_buffer_i3 (.D(quad_count[3]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i3.GSR = "DISABLED";
    FD1S3AX quad_buffer_i2 (.D(quad_count[2]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i2.GSR = "DISABLED";
    FD1S3AX quad_buffer_i1 (.D(quad_count[1]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i1.GSR = "DISABLED";
    FD1S3AX AB_i1 (.D(sync[1]), .CK(clk_1MHz), .Q(AB[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam AB_i1.GSR = "DISABLED";
    FD1S3AX sync_i1 (.D(\quad_a[2] ), .CK(clk_1MHz), .Q(sync[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam sync_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_1547[31] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i31 (.D(\spi_data_out_r_39__N_1547[30] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i30 (.D(\spi_data_out_r_39__N_1547[29] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i29 (.D(\spi_data_out_r_39__N_1547[28] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i28 (.D(\spi_data_out_r_39__N_1547[27] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i27 (.D(\spi_data_out_r_39__N_1547[26] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i26 (.D(\spi_data_out_r_39__N_1547[25] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i25 (.D(\spi_data_out_r_39__N_1547[24] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i24 (.D(\spi_data_out_r_39__N_1547[23] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i23 (.D(\spi_data_out_r_39__N_1547[22] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i22 (.D(\spi_data_out_r_39__N_1547[21] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i21 (.D(\spi_data_out_r_39__N_1547[20] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i20 (.D(\spi_data_out_r_39__N_1547[19] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i19 (.D(\spi_data_out_r_39__N_1547[18] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i18 (.D(\spi_data_out_r_39__N_1547[17] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i17 (.D(\spi_data_out_r_39__N_1547[16] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i16 (.D(\spi_data_out_r_39__N_1547[15] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_1547[14] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_1547[13] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_1547[12] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_1547[11] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_1547[10] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_1547[9] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_1547[8] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_1547[7] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_1547[6] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_1547[5] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_1547[4] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_1547[3] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_1547[2] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_1547[1] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1402[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i31 (.D(n14_adj_7176), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i31.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i30 (.D(n14_adj_7177), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i30.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i29 (.D(n14_adj_7178), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i29.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i28 (.D(n14_adj_7179), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i28.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i27 (.D(n14_adj_7180), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i27.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i26 (.D(n14_adj_7181), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i26.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i25 (.D(n14_adj_7182), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i25.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i24 (.D(n14_adj_7183), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i24.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i23 (.D(n14_adj_7184), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i23.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i22 (.D(n14_adj_7185), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i22.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i21 (.D(n14_adj_7186), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i21.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i20 (.D(n14_adj_7187), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i20.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i19 (.D(n14_adj_7188), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i19.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i18 (.D(n14_adj_7189), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i18.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i17 (.D(n14_adj_7190), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i17.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i16 (.D(n14_adj_7191), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i16.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i15 (.D(n14_adj_7192), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i15.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i14 (.D(n14_adj_7193), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i14.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i13 (.D(n14_adj_7194), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i13.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i12 (.D(n14_adj_7195), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i12.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i11 (.D(n14_adj_7196), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i11.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i10 (.D(n14_adj_7197), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i10.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i9 (.D(n14_adj_7198), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i9.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i8 (.D(n14_adj_7199), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i8.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i7 (.D(n14_adj_7200), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i7.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i6 (.D(n14_adj_7201), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i6.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i5 (.D(n14_adj_7202), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i5.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i4 (.D(n14_adj_7203), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i4.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i3 (.D(n14_adj_7204), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i3.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i2 (.D(n14_adj_7205), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i1 (.D(n14_adj_7206), .SP(clk_1MHz_enable_278), 
            .CK(clk_1MHz), .Q(quad_count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i1.GSR = "DISABLED";
    LUT4 i33_4_lut (.A(n6301[31]), .B(quad_set[31]), .C(n3_c), .D(n27301), 
         .Z(n14_adj_7176)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_907 (.A(n6301[30]), .B(quad_set[30]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7177)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_907.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_908 (.A(n6301[29]), .B(quad_set[29]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7178)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_908.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_909 (.A(n6301[28]), .B(quad_set[28]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7179)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_909.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_910 (.A(n6301[27]), .B(quad_set[27]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7180)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_910.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_911 (.A(n6301[26]), .B(quad_set[26]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7181)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_911.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_912 (.A(n6301[25]), .B(quad_set[25]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7182)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_912.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_913 (.A(n6301[24]), .B(quad_set[24]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7183)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_913.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_914 (.A(n6301[23]), .B(quad_set[23]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7184)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_914.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_915 (.A(n6301[22]), .B(quad_set[22]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7185)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_915.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_916 (.A(n6301[21]), .B(quad_set[21]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7186)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_916.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_917 (.A(n6301[20]), .B(quad_set[20]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7187)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_917.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_918 (.A(n6301[19]), .B(quad_set[19]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7188)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_918.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_919 (.A(n6301[18]), .B(quad_set[18]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7189)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_919.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_920 (.A(n6301[17]), .B(quad_set[17]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7190)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_920.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_921 (.A(n6301[16]), .B(quad_set[16]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7191)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_921.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_922 (.A(n6301[15]), .B(quad_set[15]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7192)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_922.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_923 (.A(n6301[14]), .B(quad_set[14]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7193)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_923.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_924 (.A(n6301[13]), .B(quad_set[13]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7194)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_924.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_925 (.A(n6301[12]), .B(quad_set[12]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7195)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_925.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_926 (.A(n6301[11]), .B(quad_set[11]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7196)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_926.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_927 (.A(n6301[10]), .B(quad_set[10]), .C(n3_c), 
         .D(n27301), .Z(n14_adj_7197)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_927.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_928 (.A(n6301[9]), .B(quad_set[9]), .C(n3_c), .D(n27301), 
         .Z(n14_adj_7198)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_928.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_929 (.A(n6301[8]), .B(quad_set[8]), .C(n3_c), .D(n27301), 
         .Z(n14_adj_7199)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_929.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_930 (.A(n6301[7]), .B(quad_set[7]), .C(n3_c), .D(n27301), 
         .Z(n14_adj_7200)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_930.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_931 (.A(n6301[6]), .B(quad_set[6]), .C(n3_c), .D(n27301), 
         .Z(n14_adj_7201)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_931.init = 16'hc0ca;
    FD1P3IX quad_homing__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_435), .CD(n29239), 
            .CK(clk), .Q(quad_homing[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam quad_homing__i1.GSR = "DISABLED";
    LUT4 i33_4_lut_adj_932 (.A(n6301[5]), .B(quad_set[5]), .C(n3_c), .D(n27301), 
         .Z(n14_adj_7202)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_932.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_933 (.A(n6301[4]), .B(quad_set[4]), .C(n3_c), .D(n27301), 
         .Z(n14_adj_7203)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_933.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_934 (.A(n6301[3]), .B(quad_set[3]), .C(n3_c), .D(n27301), 
         .Z(n14_adj_7204)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_934.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_935 (.A(n6301[2]), .B(quad_set[2]), .C(n3_c), .D(n27301), 
         .Z(n14_adj_7205)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_935.init = 16'hc0ca;
    LUT4 i33_4_lut_adj_936 (.A(n6301[1]), .B(quad_set[1]), .C(n3_c), .D(n27301), 
         .Z(n14_adj_7206)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_936.init = 16'hc0ca;
    FD1P3IX quad_set_valid_404 (.D(n29122), .SP(clk_enable_503), .CD(n29239), 
            .CK(clk), .Q(quad_set_valid_c)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set_valid_404.GSR = "DISABLED";
    CCU2D add_2046_33 (.A0(resetn_c), .B0(n11606), .C0(quad_count[30]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[31]), 
          .D1(GND_net), .CIN(n25150), .S0(n6301[30]), .S1(n6301[31]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_33.INIT0 = 16'hd2d2;
    defparam add_2046_33.INIT1 = 16'hd2d2;
    defparam add_2046_33.INJECT1_0 = "NO";
    defparam add_2046_33.INJECT1_1 = "NO";
    CCU2D add_2046_31 (.A0(resetn_c), .B0(n11606), .C0(quad_count[28]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[29]), 
          .D1(GND_net), .CIN(n25149), .COUT(n25150), .S0(n6301[28]), 
          .S1(n6301[29]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_31.INIT0 = 16'hd2d2;
    defparam add_2046_31.INIT1 = 16'hd2d2;
    defparam add_2046_31.INJECT1_0 = "NO";
    defparam add_2046_31.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(n29326), .B(resetn_c), .C(n108), .D(quad_set_valid), 
         .Z(n3)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/s_links/sources/mcm_top.v(17[27:33])
    defparam i2_4_lut.init = 16'h8000;
    CCU2D add_2046_29 (.A0(resetn_c), .B0(n11606), .C0(quad_count[26]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[27]), 
          .D1(GND_net), .CIN(n25148), .COUT(n25149), .S0(n6301[26]), 
          .S1(n6301[27]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_29.INIT0 = 16'hd2d2;
    defparam add_2046_29.INIT1 = 16'hd2d2;
    defparam add_2046_29.INJECT1_0 = "NO";
    defparam add_2046_29.INJECT1_1 = "NO";
    CCU2D add_2046_27 (.A0(resetn_c), .B0(n11606), .C0(quad_count[24]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[25]), 
          .D1(GND_net), .CIN(n25147), .COUT(n25148), .S0(n6301[24]), 
          .S1(n6301[25]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_27.INIT0 = 16'hd2d2;
    defparam add_2046_27.INIT1 = 16'hd2d2;
    defparam add_2046_27.INJECT1_0 = "NO";
    defparam add_2046_27.INJECT1_1 = "NO";
    CCU2D add_2046_25 (.A0(resetn_c), .B0(n11606), .C0(quad_count[22]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[23]), 
          .D1(GND_net), .CIN(n25146), .COUT(n25147), .S0(n6301[22]), 
          .S1(n6301[23]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_25.INIT0 = 16'hd2d2;
    defparam add_2046_25.INIT1 = 16'hd2d2;
    defparam add_2046_25.INJECT1_0 = "NO";
    defparam add_2046_25.INJECT1_1 = "NO";
    CCU2D add_2046_23 (.A0(resetn_c), .B0(n11606), .C0(quad_count[20]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[21]), 
          .D1(GND_net), .CIN(n25145), .COUT(n25146), .S0(n6301[20]), 
          .S1(n6301[21]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_23.INIT0 = 16'hd2d2;
    defparam add_2046_23.INIT1 = 16'hd2d2;
    defparam add_2046_23.INJECT1_0 = "NO";
    defparam add_2046_23.INJECT1_1 = "NO";
    CCU2D add_2046_21 (.A0(resetn_c), .B0(n11606), .C0(quad_count[18]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[19]), 
          .D1(GND_net), .CIN(n25144), .COUT(n25145), .S0(n6301[18]), 
          .S1(n6301[19]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_21.INIT0 = 16'hd2d2;
    defparam add_2046_21.INIT1 = 16'hd2d2;
    defparam add_2046_21.INJECT1_0 = "NO";
    defparam add_2046_21.INJECT1_1 = "NO";
    CCU2D add_2046_19 (.A0(resetn_c), .B0(n11606), .C0(quad_count[16]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[17]), 
          .D1(GND_net), .CIN(n25143), .COUT(n25144), .S0(n6301[16]), 
          .S1(n6301[17]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_19.INIT0 = 16'hd2d2;
    defparam add_2046_19.INIT1 = 16'hd2d2;
    defparam add_2046_19.INJECT1_0 = "NO";
    defparam add_2046_19.INJECT1_1 = "NO";
    CCU2D add_2046_17 (.A0(resetn_c), .B0(n11606), .C0(quad_count[14]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[15]), 
          .D1(GND_net), .CIN(n25142), .COUT(n25143), .S0(n6301[14]), 
          .S1(n6301[15]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_17.INIT0 = 16'hd2d2;
    defparam add_2046_17.INIT1 = 16'hd2d2;
    defparam add_2046_17.INJECT1_0 = "NO";
    defparam add_2046_17.INJECT1_1 = "NO";
    CCU2D add_2046_15 (.A0(resetn_c), .B0(n11606), .C0(quad_count[12]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[13]), 
          .D1(GND_net), .CIN(n25141), .COUT(n25142), .S0(n6301[12]), 
          .S1(n6301[13]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_15.INIT0 = 16'hd2d2;
    defparam add_2046_15.INIT1 = 16'hd2d2;
    defparam add_2046_15.INJECT1_0 = "NO";
    defparam add_2046_15.INJECT1_1 = "NO";
    CCU2D add_2046_13 (.A0(resetn_c), .B0(n11606), .C0(quad_count[10]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[11]), 
          .D1(GND_net), .CIN(n25140), .COUT(n25141), .S0(n6301[10]), 
          .S1(n6301[11]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_13.INIT0 = 16'hd2d2;
    defparam add_2046_13.INIT1 = 16'hd2d2;
    defparam add_2046_13.INJECT1_0 = "NO";
    defparam add_2046_13.INJECT1_1 = "NO";
    CCU2D add_2046_11 (.A0(resetn_c), .B0(n11606), .C0(quad_count[8]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[9]), 
          .D1(GND_net), .CIN(n25139), .COUT(n25140), .S0(n6301[8]), 
          .S1(n6301[9]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_11.INIT0 = 16'hd2d2;
    defparam add_2046_11.INIT1 = 16'hd2d2;
    defparam add_2046_11.INJECT1_0 = "NO";
    defparam add_2046_11.INJECT1_1 = "NO";
    CCU2D add_2046_9 (.A0(resetn_c), .B0(n11606), .C0(quad_count[6]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[7]), 
          .D1(GND_net), .CIN(n25138), .COUT(n25139), .S0(n6301[6]), 
          .S1(n6301[7]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_9.INIT0 = 16'hd2d2;
    defparam add_2046_9.INIT1 = 16'hd2d2;
    defparam add_2046_9.INJECT1_0 = "NO";
    defparam add_2046_9.INJECT1_1 = "NO";
    CCU2D add_2046_7 (.A0(resetn_c), .B0(n11606), .C0(quad_count[4]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[5]), 
          .D1(GND_net), .CIN(n25137), .COUT(n25138), .S0(n6301[4]), 
          .S1(n6301[5]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_7.INIT0 = 16'hd2d2;
    defparam add_2046_7.INIT1 = 16'hd2d2;
    defparam add_2046_7.INJECT1_0 = "NO";
    defparam add_2046_7.INJECT1_1 = "NO";
    CCU2D add_2046_5 (.A0(resetn_c), .B0(n11606), .C0(quad_count[2]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[3]), 
          .D1(GND_net), .CIN(n25136), .COUT(n25137), .S0(n6301[2]), 
          .S1(n6301[3]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_5.INIT0 = 16'hd2d2;
    defparam add_2046_5.INIT1 = 16'hd2d2;
    defparam add_2046_5.INJECT1_0 = "NO";
    defparam add_2046_5.INJECT1_1 = "NO";
    CCU2D add_2046_3 (.A0(resetn_c), .B0(n11606), .C0(quad_count[0]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11606), .C1(quad_count[1]), 
          .D1(GND_net), .CIN(n25135), .COUT(n25136), .S0(n6301[0]), 
          .S1(n6301[1]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_3.INIT0 = 16'h2d2d;
    defparam add_2046_3.INIT1 = 16'hd2d2;
    defparam add_2046_3.INJECT1_0 = "NO";
    defparam add_2046_3.INJECT1_1 = "NO";
    CCU2D add_2046_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(resetn_c), .B1(n11606), .C1(GND_net), .D1(GND_net), .COUT(n25135));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2046_1.INIT0 = 16'hF000;
    defparam add_2046_1.INIT1 = 16'hdddd;
    defparam add_2046_1.INJECT1_0 = "NO";
    defparam add_2046_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(resetn_c), .B(mem_rdata_update_N_729), .Z(n9633)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/mcm_top.v(17[27:33])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i22915_4_lut (.A(resetn_c), .B(n12714), .C(n26751), .D(quad_set_valid_c), 
         .Z(clk_1MHz_enable_278)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i22915_4_lut.init = 16'hffdf;
    LUT4 i33_4_lut_adj_937 (.A(n6301[0]), .B(quad_set[0]), .C(n3_c), .D(n27301), 
         .Z(n14)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_937.init = 16'hc0ca;
    LUT4 i1_4_lut (.A(quad_set_valid_c), .B(n36), .C(n13), .D(n29053), 
         .Z(n3_c)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_4_lut.init = 16'h8880;
    LUT4 i2_4_lut_adj_938 (.A(n12820), .B(n1711[2]), .C(n1711[1]), .D(n29234), 
         .Z(n13)) /* synthesis lut_function=(!((B+!(C (D)+!C !(D)))+!A)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i2_4_lut_adj_938.init = 16'h2002;
    LUT4 i1_2_lut_adj_939 (.A(resetn_c), .B(n1711[3]), .Z(n12820)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_939.init = 16'h2222;
    LUT4 i1_2_lut_adj_940 (.A(n1711[2]), .B(n1711[1]), .Z(n59)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i1_2_lut_adj_940.init = 16'heeee;
    LUT4 i1_2_lut_adj_941 (.A(n1711[0]), .B(n1711[3]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam i1_2_lut_adj_941.init = 16'heeee;
    LUT4 n59_bdd_4_lut (.A(n59), .B(n1711[0]), .C(AB[1]), .D(AB[0]), 
         .Z(n28870)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D)))) */ ;
    defparam n59_bdd_4_lut.init = 16'hc00e;
    LUT4 i2_4_lut_adj_942 (.A(n29336), .B(resetn_c), .C(n95), .D(quad_set_valid_adj_207), 
         .Z(n5647)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/s_links/sources/mcm_top.v(17[27:33])
    defparam i2_4_lut_adj_942.init = 16'h8000;
    
endmodule
//
// Verilog Description of module pll
//

module pll (clk_in_c, clk_1MHz, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input clk_in_c;
    output clk_1MHz;
    input GND_net;
    
    wire clk_in_c /* synthesis is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(16[27:33])
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    
    wire CLKFB_t;
    
    EHXPLLJ PLLInst_0 (.CLKI(clk_in_c), .CLKFB(CLKFB_t), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(GND_net), .PLLRST(GND_net), .PLLSTB(GND_net), 
            .PLLWE(GND_net), .PLLDATI0(GND_net), .PLLDATI1(GND_net), .PLLDATI2(GND_net), 
            .PLLDATI3(GND_net), .PLLDATI4(GND_net), .PLLDATI5(GND_net), 
            .PLLDATI6(GND_net), .PLLDATI7(GND_net), .PLLADDR0(GND_net), 
            .PLLADDR1(GND_net), .PLLADDR2(GND_net), .PLLADDR3(GND_net), 
            .PLLADDR4(GND_net), .CLKOS3(clk_1MHz), .CLKINTFB(CLKFB_t)) /* synthesis FREQUENCY_PIN_CLKOS3="1.000000", FREQUENCY_PIN_CLKOS2="0.020000", FREQUENCY_PIN_CLKOS="0.100000", FREQUENCY_PIN_CLKOP="96.000000", FREQUENCY_PIN_CLKI="12.000000", ICP_CURRENT="9", LPF_RESISTOR="4", syn_instantiated=1, LSE_LINE_FILE_ID=3, LSE_LCOL=5, LSE_RCOL=100, LSE_LLINE=149, LSE_RLINE=149 */ ;   // c:/s_links/sources/mcm_top.v(149[5:100])
    defparam PLLInst_0.CLKI_DIV = 1;
    defparam PLLInst_0.CLKFB_DIV = 8;
    defparam PLLInst_0.CLKOP_DIV = 3;
    defparam PLLInst_0.CLKOS_DIV = 120;
    defparam PLLInst_0.CLKOS2_DIV = 120;
    defparam PLLInst_0.CLKOS3_DIV = 12;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "ENABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "ENABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "ENABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 2;
    defparam PLLInst_0.CLKOS_CPHASE = 119;
    defparam PLLInst_0.CLKOS2_CPHASE = 119;
    defparam PLLInst_0.CLKOS3_CPHASE = 11;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "INT_DIVA";
    defparam PLLInst_0.FRACN_ENABLE = "DISABLED";
    defparam PLLInst_0.FRACN_DIV = 0;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "DISABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 3;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module \piezo(DEV_ID=6,UART_ADDRESS_WIDTH=4) 
//

module \piezo(DEV_ID=6,UART_ADDRESS_WIDTH=4)  (n28811, n28813, mode, clk, 
            clk_enable_188, n29239, n29762, n29191, n29190, pin_io_out_65, 
            n25382, pin_io_out_26, pin_io_out_16, n29157, n7, pin_io_out_40, 
            n29189, C_8_c, tx_N_6443, pin_io_out_45, n27189, pin_io_out_46, 
            pin_io_out_55, n29150, n27186, n29202, pin_io_out_15, 
            n29198, n13, pin_io_out_56, n29196, n29158, n26972, 
            n22, pin_io_out_5, n29160, n29153, n26951, n14, OW_ID_N_4464, 
            n27480, n27483, n29132, n27471, n29199, n27477, mode_adj_183, 
            mode_adj_184, n29203, mode_adj_185, mode_adj_186, C_2_c_1, 
            C_1_c_0, C_5_c_c, n29313, mode_adj_187, n29284, mode_adj_188, 
            mode_adj_189, mode_adj_190, pin_io_out_25, n22_adj_191, 
            mode_adj_192, mode_adj_193, n31, mode_adj_194, mode_adj_195, 
            n29285, \cs_decoded[8] , n5, mode_adj_196, n29293, mode_adj_197, 
            mode_adj_198, n29299, n29301, \mode[0] , n8679, n29305, 
            \mode[1] , n29300, n29317, n8739, \cs_decoded[6] , n8740, 
            mode_adj_199, mode_adj_200, n29303, \cs_decoded[4] , n29295, 
            n8768, \cs_decoded[13] , n2, n8836, mode_adj_206, digital_output_r, 
            n26521, n29267, mode_adj_203, pin_io_out_66, mode_adj_204, 
            pin_io_out_36, mode_adj_205) /* synthesis syn_module_defined=1 */ ;
    input n28811;
    output n28813;
    output mode;
    input clk;
    input clk_enable_188;
    input n29239;
    input n29762;
    input n29191;
    input n29190;
    input pin_io_out_65;
    output n25382;
    input pin_io_out_26;
    input pin_io_out_16;
    input n29157;
    input n7;
    input pin_io_out_40;
    input n29189;
    input C_8_c;
    input tx_N_6443;
    input pin_io_out_45;
    input n27189;
    input pin_io_out_46;
    input pin_io_out_55;
    input n29150;
    input n27186;
    input n29202;
    input pin_io_out_15;
    input n29198;
    output n13;
    input pin_io_out_56;
    input n29196;
    input n29158;
    input n26972;
    input n22;
    input pin_io_out_5;
    input n29160;
    input n29153;
    output n26951;
    input n14;
    input OW_ID_N_4464;
    input n27480;
    input n27483;
    input n29132;
    input n27471;
    input n29199;
    input n27477;
    input mode_adj_183;
    input mode_adj_184;
    input n29203;
    input mode_adj_185;
    input mode_adj_186;
    input C_2_c_1;
    input C_1_c_0;
    input C_5_c_c;
    input n29313;
    input mode_adj_187;
    input n29284;
    input mode_adj_188;
    input mode_adj_189;
    input mode_adj_190;
    input pin_io_out_25;
    input n22_adj_191;
    input mode_adj_192;
    input mode_adj_193;
    output n31;
    input mode_adj_194;
    input mode_adj_195;
    output n29285;
    input \cs_decoded[8] ;
    output n5;
    input mode_adj_196;
    output n29293;
    input mode_adj_197;
    input mode_adj_198;
    output n29299;
    input n29301;
    input \mode[0] ;
    output n8679;
    input n29305;
    input \mode[1] ;
    output n29300;
    input n29317;
    output n8739;
    input \cs_decoded[6] ;
    output n8740;
    input mode_adj_199;
    input mode_adj_200;
    output n29303;
    input \cs_decoded[4] ;
    input n29295;
    output n8768;
    input \cs_decoded[13] ;
    output n2;
    output n8836;
    input [2:0]mode_adj_206;
    input digital_output_r;
    output n26521;
    input n29267;
    input mode_adj_203;
    input pin_io_out_66;
    input mode_adj_204;
    input pin_io_out_36;
    input mode_adj_205;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    wire n28812, n19229, n34, n17, n30, n26, n29335, n29151, 
        n27, n28, n22_c, n20, n25329, n26977, n24, n27950, n18, 
        n20_adj_7152, n10, n8, n27467, n32, n29276, n29334, n29333;
    
    PFUMX i23079 (.BLUT(n28812), .ALUT(n28811), .C0(n19229), .Z(n28813));
    FD1P3IX mode_38 (.D(n29762), .SP(clk_enable_188), .CD(n29239), .CK(clk), 
            .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=632, LSE_RLINE=661 */ ;   // c:/s_links/sources/slot_cards/piezo.v(55[8] 63[4])
    defparam mode_38.GSR = "DISABLED";
    LUT4 Select_3812_i34_2_lut_4_lut (.A(n29191), .B(n29190), .C(mode), 
         .D(pin_io_out_65), .Z(n34)) /* synthesis lut_function=(!(A+!(B (D)+!B (C (D))))) */ ;   // c:/s_links/sources/slot_cards/piezo.v(51[8:15])
    defparam Select_3812_i34_2_lut_4_lut.init = 16'h5400;
    LUT4 i15_4_lut (.A(n17), .B(n30), .C(n26), .D(n29335), .Z(n25382)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut (.A(pin_io_out_26), .B(pin_io_out_16), .C(n29151), .D(n29157), 
         .Z(n17)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i14_4_lut (.A(n27), .B(n28), .C(n22_c), .D(n7), .Z(n30)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i10_4_lut (.A(pin_io_out_40), .B(n20), .C(n25329), .D(n29189), 
         .Z(n26)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut.init = 16'hfefc;
    LUT4 Select_3812_i27_2_lut (.A(C_8_c), .B(tx_N_6443), .Z(n27)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam Select_3812_i27_2_lut.init = 16'h2222;
    LUT4 i12_4_lut (.A(n26977), .B(n24), .C(pin_io_out_45), .D(n27189), 
         .Z(n28)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i12_4_lut.init = 16'hfeee;
    LUT4 i6_4_lut (.A(pin_io_out_46), .B(pin_io_out_55), .C(n29150), .D(n27186), 
         .Z(n22_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut.init = 16'heca0;
    LUT4 i1_4_lut_adj_902 (.A(n29202), .B(pin_io_out_15), .C(n29198), 
         .D(n13), .Z(n26977)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;
    defparam i1_4_lut_adj_902.init = 16'h4440;
    LUT4 i8_4_lut (.A(pin_io_out_56), .B(n29196), .C(n29158), .D(n26972), 
         .Z(n24)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A !(B+!(D))) */ ;
    defparam i8_4_lut.init = 16'hb3a0;
    LUT4 i4_4_lut (.A(n22), .B(n34), .C(pin_io_out_5), .D(n29160), .Z(n20)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i4_4_lut.init = 16'hccec;
    LUT4 i22791_4_lut (.A(n29153), .B(n27950), .C(n18), .D(tx_N_6443), 
         .Z(n26951)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i22791_4_lut.init = 16'h0400;
    LUT4 i22790_4_lut (.A(n29158), .B(n20_adj_7152), .C(n14), .D(n29157), 
         .Z(n27950)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i22790_4_lut.init = 16'h0001;
    LUT4 i6_4_lut_adj_903 (.A(OW_ID_N_4464), .B(n27480), .C(n10), .D(n27483), 
         .Z(n18)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut_adj_903.init = 16'hfffe;
    LUT4 i8_4_lut_adj_904 (.A(n29151), .B(n29189), .C(n29132), .D(n29150), 
         .Z(n20_adj_7152)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i8_4_lut_adj_904.init = 16'hfffe;
    LUT4 i4_4_lut_adj_905 (.A(n29196), .B(n8), .C(n27471), .D(n27467), 
         .Z(n10)) /* synthesis lut_function=(A (B+(C))+!A (B+(C+(D)))) */ ;
    defparam i4_4_lut_adj_905.init = 16'hfdfc;
    LUT4 i2_4_lut (.A(n29199), .B(n27477), .C(mode_adj_183), .D(n32), 
         .Z(n8)) /* synthesis lut_function=(A (B)+!A (B+(C+(D)))) */ ;
    defparam i2_4_lut.init = 16'hdddc;
    LUT4 i22_4_lut (.A(mode_adj_184), .B(n29203), .C(mode_adj_185), .D(mode_adj_186), 
         .Z(n27467)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_548 (.A(C_2_c_1), .B(C_1_c_0), .Z(n29276)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam i1_2_lut_rep_548.init = 16'hbbbb;
    LUT4 i14302_2_lut_3_lut_4_lut (.A(C_2_c_1), .B(C_1_c_0), .C(C_5_c_c), 
         .D(n29313), .Z(n19229)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam i14302_2_lut_3_lut_4_lut.init = 16'hfbff;
    LUT4 OW_ID_I_263_2_lut_rep_423_3_lut_4_lut (.A(C_2_c_1), .B(C_1_c_0), 
         .C(mode_adj_187), .D(n29284), .Z(n29151)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam OW_ID_I_263_2_lut_rep_423_3_lut_4_lut.init = 16'h0040;
    LUT4 i5_3_lut (.A(mode_adj_188), .B(mode_adj_189), .C(mode_adj_190), 
         .Z(n13)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i5_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_4_lut (.A(n29284), .B(n29276), .C(pin_io_out_25), .D(n22_adj_191), 
         .Z(n25329)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/s_links/sources/slot_cards/piezo.v(50[44:72])
    defparam i2_3_lut_4_lut.init = 16'h1000;
    LUT4 i11_2_lut (.A(mode_adj_192), .B(mode_adj_193), .Z(n31)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i11_2_lut.init = 16'heeee;
    LUT4 i12_2_lut_rep_557 (.A(mode_adj_194), .B(mode_adj_195), .Z(n29285)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12_2_lut_rep_557.init = 16'heeee;
    LUT4 Select_3926_i5_2_lut_3_lut (.A(mode_adj_194), .B(mode_adj_195), 
         .C(\cs_decoded[8] ), .Z(n5)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam Select_3926_i5_2_lut_3_lut.init = 16'he0e0;
    LUT4 i3870_2_lut_rep_565 (.A(mode_adj_196), .B(mode), .Z(n29293)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/piezo.v(46[8:14])
    defparam i3870_2_lut_rep_565.init = 16'heeee;
    LUT4 i7_2_lut_rep_571 (.A(mode_adj_197), .B(mode_adj_198), .Z(n29299)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7_2_lut_rep_571.init = 16'heeee;
    LUT4 i22759_2_lut_2_lut_3_lut_4_lut (.A(mode_adj_197), .B(mode_adj_198), 
         .C(n29301), .D(\mode[0] ), .Z(n8679)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;
    defparam i22759_2_lut_2_lut_3_lut_4_lut.init = 16'h1011;
    LUT4 i15_2_lut_3_lut_4_lut (.A(mode_adj_197), .B(mode_adj_198), .C(n29305), 
         .D(\mode[1] ), .Z(n32)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i15_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i13_2_lut_rep_572 (.A(mode_adj_185), .B(mode_adj_186), .Z(n29300)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13_2_lut_rep_572.init = 16'heeee;
    LUT4 i22735_2_lut_2_lut_3_lut (.A(mode_adj_185), .B(mode_adj_186), .C(n29317), 
         .Z(n8739)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i22735_2_lut_2_lut_3_lut.init = 16'h0101;
    LUT4 Select_3958_i7_3_lut_4_lut (.A(mode_adj_185), .B(mode_adj_186), 
         .C(\cs_decoded[6] ), .D(n29317), .Z(n8740)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;
    defparam Select_3958_i7_3_lut_4_lut.init = 16'hffe0;
    LUT4 i2_2_lut_rep_575 (.A(mode_adj_199), .B(mode_adj_200), .Z(n29303)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut_rep_575.init = 16'heeee;
    LUT4 Select_3986_i7_3_lut_4_lut (.A(mode_adj_199), .B(mode_adj_200), 
         .C(\cs_decoded[4] ), .D(n29295), .Z(n8768)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(D))) */ ;
    defparam Select_3986_i7_3_lut_4_lut.init = 16'he0ff;
    LUT4 Select_3863_i2_2_lut (.A(\cs_decoded[13] ), .B(mode), .Z(n2)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_3863_i2_2_lut.init = 16'h8888;
    LUT4 i4121_1_lut (.A(mode), .Z(n8836)) /* synthesis lut_function=(!(A)) */ ;
    defparam i4121_1_lut.init = 16'h5555;
    LUT4 i3_4_lut (.A(mode_adj_206[2]), .B(digital_output_r), .C(mode_adj_206[1]), 
         .D(mode_adj_206[0]), .Z(n26521)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i3_4_lut.init = 16'h4000;
    LUT4 RESET_N_6154_bdd_4_lut (.A(n29267), .B(mode_adj_203), .C(n29293), 
         .D(mode_adj_206[0]), .Z(n28812)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam RESET_N_6154_bdd_4_lut.init = 16'h0002;
    LUT4 i2_4_lut_then_4_lut (.A(pin_io_out_66), .B(C_2_c_1), .C(n29313), 
         .D(mode_adj_204), .Z(n29334)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i2_4_lut_then_4_lut.init = 16'h2000;
    LUT4 i2_4_lut_else_4_lut (.A(pin_io_out_36), .B(C_2_c_1), .C(n29284), 
         .D(mode_adj_205), .Z(n29333)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2_4_lut_else_4_lut.init = 16'h0800;
    PFUMX i23164 (.BLUT(n29333), .ALUT(n29334), .C0(C_1_c_0), .Z(n29335));
    
endmodule
//
// Verilog Description of module \intrpt_ctrl(DEV_ID=6) 
//

module \intrpt_ctrl(DEV_ID=6)  (clk, n29239, \spi_data_out_r_39__N_2998[0] , 
            \pin_intrpt[18] , \pin_intrpt[20] , \pin_intrpt[19] , clear_intrpt, 
            clear_intrpt_N_3065, intrpt_out_c_6, intrpt_out_N_3061, n29757, 
            \spi_data_out_r_39__N_2998[2] , \spi_data_out_r_39__N_2998[1] ) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input n29239;
    output \spi_data_out_r_39__N_2998[0] ;
    input \pin_intrpt[18] ;
    input \pin_intrpt[20] ;
    input \pin_intrpt[19] ;
    output clear_intrpt;
    input clear_intrpt_N_3065;
    output intrpt_out_c_6;
    input intrpt_out_N_3061;
    input n29757;
    output \spi_data_out_r_39__N_2998[2] ;
    output \spi_data_out_r_39__N_2998[1] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire \pin_intrpt[20]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[20] */ ;   // c:/s_links/sources/mcm_top.v(102[46:56])
    wire [2:0]intrpt_in_dly;   // c:/s_links/sources/intrpt_ctrl.v(39[36:49])
    wire [2:0]intrpt_in_reg;   // c:/s_links/sources/intrpt_ctrl.v(38[35:48])
    
    wire assert_intrpt, intrpt_all_edges, n4;
    
    FD1S3IX intrpt_in_dly__i0 (.D(intrpt_in_reg[0]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\pin_intrpt[18] ), .CK(clk), .Q(\spi_data_out_r_39__N_2998[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i0 (.D(\pin_intrpt[18] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i0.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i2 (.D(\pin_intrpt[20] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_reg__i1 (.D(\pin_intrpt[19] ), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_reg[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(49[8] 54[4])
    defparam intrpt_in_reg__i1.GSR = "DISABLED";
    FD1S3IX clear_intrpt_317 (.D(clear_intrpt_N_3065), .CK(clk), .CD(n29239), 
            .Q(clear_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam clear_intrpt_317.GSR = "DISABLED";
    FD1S3IX assert_intrpt_316 (.D(intrpt_all_edges), .CK(clk), .CD(n29239), 
            .Q(assert_intrpt)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(63[8] 73[4])
    defparam assert_intrpt_316.GSR = "DISABLED";
    FD1P3IX intrpt_out_359 (.D(n29757), .SP(assert_intrpt), .CD(intrpt_out_N_3061), 
            .CK(clk), .Q(intrpt_out_c_6)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(92[8] 99[4])
    defparam intrpt_out_359.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\pin_intrpt[20] ), .CK(clk), .Q(\spi_data_out_r_39__N_2998[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\pin_intrpt[19] ), .CK(clk), .Q(\spi_data_out_r_39__N_2998[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(78[8] 89[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i2 (.D(intrpt_in_reg[2]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i2.GSR = "DISABLED";
    FD1S3IX intrpt_in_dly__i1 (.D(intrpt_in_reg[1]), .CK(clk), .CD(n29239), 
            .Q(intrpt_in_dly[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=304, LSE_RLINE=325 */ ;   // c:/s_links/sources/intrpt_ctrl.v(56[8] 61[4])
    defparam intrpt_in_dly__i1.GSR = "DISABLED";
    LUT4 i2_3_lut (.A(intrpt_in_dly[0]), .B(n4), .C(intrpt_in_reg[0]), 
         .Z(intrpt_all_edges)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i2_3_lut.init = 16'hdede;
    LUT4 i1_4_lut (.A(intrpt_in_dly[1]), .B(intrpt_in_dly[2]), .C(intrpt_in_reg[1]), 
         .D(intrpt_in_reg[2]), .Z(n4)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;   // c:/s_links/sources/intrpt_ctrl.v(47[27:74])
    defparam i1_4_lut.init = 16'h7bde;
    
endmodule
//
// Verilog Description of module \quad_decoder(DEV_ID=3) 
//

module \quad_decoder(DEV_ID=3)  (quad_count, clk_1MHz, \spi_data_out_r_39__N_1636[0] , 
            clk, \spi_data_out_r_39__N_1781[0] , \quad_b[3] , quad_buffer, 
            \pin_intrpt[11] , clk_enable_398, n29239, \spi_data_r[0] , 
            clk_enable_434, n29762, quad_set_complete, spi_data_out_r_39__N_1676, 
            n29098, \spi_addr[0] , n26933, n13511, spi_data_out_r_39__N_2332, 
            n13506, spi_data_out_r_39__N_1396, n13413, \quad_a[3] , 
            \spi_data_out_r_39__N_1636[31] , \spi_data_out_r_39__N_1781[31] , 
            resetn_c, GND_net, \spi_data_out_r_39__N_1636[30] , \spi_data_out_r_39__N_1781[30] , 
            \spi_data_out_r_39__N_1636[29] , \spi_data_out_r_39__N_1781[29] , 
            \spi_data_out_r_39__N_1636[28] , \spi_data_out_r_39__N_1781[28] , 
            \spi_data_out_r_39__N_1636[27] , \spi_data_out_r_39__N_1781[27] , 
            \spi_data_out_r_39__N_1636[26] , \spi_data_out_r_39__N_1781[26] , 
            \spi_data_out_r_39__N_1636[25] , \spi_data_out_r_39__N_1781[25] , 
            \spi_data_out_r_39__N_1636[24] , \spi_data_out_r_39__N_1781[24] , 
            \spi_data_out_r_39__N_1636[23] , \spi_data_out_r_39__N_1781[23] , 
            \spi_data_out_r_39__N_1636[22] , \spi_data_out_r_39__N_1781[22] , 
            \spi_data_out_r_39__N_1636[21] , \spi_data_out_r_39__N_1781[21] , 
            \spi_data_out_r_39__N_1636[20] , \spi_data_out_r_39__N_1781[20] , 
            \spi_data_out_r_39__N_1636[19] , \spi_data_out_r_39__N_1781[19] , 
            \spi_data_out_r_39__N_1636[18] , \spi_data_out_r_39__N_1781[18] , 
            \spi_data_out_r_39__N_1636[17] , \spi_data_out_r_39__N_1781[17] , 
            \spi_data_out_r_39__N_1636[16] , \spi_data_out_r_39__N_1781[16] , 
            \spi_data_out_r_39__N_1636[15] , \spi_data_out_r_39__N_1781[15] , 
            \spi_data_out_r_39__N_1636[14] , \spi_data_out_r_39__N_1781[14] , 
            \spi_data_out_r_39__N_1636[13] , \spi_data_out_r_39__N_1781[13] , 
            \spi_data_out_r_39__N_1636[12] , \spi_data_out_r_39__N_1781[12] , 
            \spi_data_out_r_39__N_1636[11] , \spi_data_out_r_39__N_1781[11] , 
            \spi_data_out_r_39__N_1636[10] , \spi_data_out_r_39__N_1781[10] , 
            \spi_data_out_r_39__N_1636[9] , \spi_data_out_r_39__N_1781[9] , 
            \spi_data_out_r_39__N_1636[8] , \spi_data_out_r_39__N_1781[8] , 
            \spi_data_out_r_39__N_1636[7] , \spi_data_out_r_39__N_1781[7] , 
            \spi_data_out_r_39__N_1636[6] , \spi_data_out_r_39__N_1781[6] , 
            \spi_data_out_r_39__N_1636[5] , \spi_data_out_r_39__N_1781[5] , 
            \spi_data_out_r_39__N_1636[4] , \spi_data_out_r_39__N_1781[4] , 
            \spi_data_out_r_39__N_1636[3] , \spi_data_out_r_39__N_1781[3] , 
            \spi_data_out_r_39__N_1636[2] , \spi_data_out_r_39__N_1781[2] , 
            \spi_data_out_r_39__N_1636[1] , \spi_data_out_r_39__N_1781[1] , 
            \spi_data_r[1] , \spi_data_r[2] , \spi_data_r[3] , \spi_data_r[4] , 
            \spi_data_r[5] , \spi_data_r[6] , \spi_data_r[7] , \spi_data_r[8] , 
            \spi_data_r[9] , \spi_data_r[10] , \spi_data_r[11] , \spi_data_r[12] , 
            \spi_data_r[13] , \spi_data_r[14] , \spi_data_r[15] , \spi_data_r[16] , 
            \spi_data_r[17] , \spi_data_r[18] , \spi_data_r[19] , \spi_data_r[20] , 
            \spi_data_r[21] , \spi_data_r[22] , \spi_data_r[23] , \spi_data_r[24] , 
            \spi_data_r[25] , \spi_data_r[26] , \spi_data_r[27] , \spi_data_r[28] , 
            \spi_data_r[29] , \spi_data_r[30] , \spi_data_r[31] , \quad_homing[1] , 
            clk_enable_505, n29120, n13052, n26969, pin_io_out_34, 
            n27632) /* synthesis syn_module_defined=1 */ ;
    output [31:0]quad_count;
    input clk_1MHz;
    output \spi_data_out_r_39__N_1636[0] ;
    input clk;
    input \spi_data_out_r_39__N_1781[0] ;
    input \quad_b[3] ;
    output [31:0]quad_buffer;
    input \pin_intrpt[11] ;
    input clk_enable_398;
    input n29239;
    input \spi_data_r[0] ;
    input clk_enable_434;
    input n29762;
    output quad_set_complete;
    output spi_data_out_r_39__N_1676;
    input n29098;
    input \spi_addr[0] ;
    input n26933;
    input n13511;
    output spi_data_out_r_39__N_2332;
    input n13506;
    output spi_data_out_r_39__N_1396;
    input n13413;
    input \quad_a[3] ;
    output \spi_data_out_r_39__N_1636[31] ;
    input \spi_data_out_r_39__N_1781[31] ;
    input resetn_c;
    input GND_net;
    output \spi_data_out_r_39__N_1636[30] ;
    input \spi_data_out_r_39__N_1781[30] ;
    output \spi_data_out_r_39__N_1636[29] ;
    input \spi_data_out_r_39__N_1781[29] ;
    output \spi_data_out_r_39__N_1636[28] ;
    input \spi_data_out_r_39__N_1781[28] ;
    output \spi_data_out_r_39__N_1636[27] ;
    input \spi_data_out_r_39__N_1781[27] ;
    output \spi_data_out_r_39__N_1636[26] ;
    input \spi_data_out_r_39__N_1781[26] ;
    output \spi_data_out_r_39__N_1636[25] ;
    input \spi_data_out_r_39__N_1781[25] ;
    output \spi_data_out_r_39__N_1636[24] ;
    input \spi_data_out_r_39__N_1781[24] ;
    output \spi_data_out_r_39__N_1636[23] ;
    input \spi_data_out_r_39__N_1781[23] ;
    output \spi_data_out_r_39__N_1636[22] ;
    input \spi_data_out_r_39__N_1781[22] ;
    output \spi_data_out_r_39__N_1636[21] ;
    input \spi_data_out_r_39__N_1781[21] ;
    output \spi_data_out_r_39__N_1636[20] ;
    input \spi_data_out_r_39__N_1781[20] ;
    output \spi_data_out_r_39__N_1636[19] ;
    input \spi_data_out_r_39__N_1781[19] ;
    output \spi_data_out_r_39__N_1636[18] ;
    input \spi_data_out_r_39__N_1781[18] ;
    output \spi_data_out_r_39__N_1636[17] ;
    input \spi_data_out_r_39__N_1781[17] ;
    output \spi_data_out_r_39__N_1636[16] ;
    input \spi_data_out_r_39__N_1781[16] ;
    output \spi_data_out_r_39__N_1636[15] ;
    input \spi_data_out_r_39__N_1781[15] ;
    output \spi_data_out_r_39__N_1636[14] ;
    input \spi_data_out_r_39__N_1781[14] ;
    output \spi_data_out_r_39__N_1636[13] ;
    input \spi_data_out_r_39__N_1781[13] ;
    output \spi_data_out_r_39__N_1636[12] ;
    input \spi_data_out_r_39__N_1781[12] ;
    output \spi_data_out_r_39__N_1636[11] ;
    input \spi_data_out_r_39__N_1781[11] ;
    output \spi_data_out_r_39__N_1636[10] ;
    input \spi_data_out_r_39__N_1781[10] ;
    output \spi_data_out_r_39__N_1636[9] ;
    input \spi_data_out_r_39__N_1781[9] ;
    output \spi_data_out_r_39__N_1636[8] ;
    input \spi_data_out_r_39__N_1781[8] ;
    output \spi_data_out_r_39__N_1636[7] ;
    input \spi_data_out_r_39__N_1781[7] ;
    output \spi_data_out_r_39__N_1636[6] ;
    input \spi_data_out_r_39__N_1781[6] ;
    output \spi_data_out_r_39__N_1636[5] ;
    input \spi_data_out_r_39__N_1781[5] ;
    output \spi_data_out_r_39__N_1636[4] ;
    input \spi_data_out_r_39__N_1781[4] ;
    output \spi_data_out_r_39__N_1636[3] ;
    input \spi_data_out_r_39__N_1781[3] ;
    output \spi_data_out_r_39__N_1636[2] ;
    input \spi_data_out_r_39__N_1781[2] ;
    output \spi_data_out_r_39__N_1636[1] ;
    input \spi_data_out_r_39__N_1781[1] ;
    input \spi_data_r[1] ;
    input \spi_data_r[2] ;
    input \spi_data_r[3] ;
    input \spi_data_r[4] ;
    input \spi_data_r[5] ;
    input \spi_data_r[6] ;
    input \spi_data_r[7] ;
    input \spi_data_r[8] ;
    input \spi_data_r[9] ;
    input \spi_data_r[10] ;
    input \spi_data_r[11] ;
    input \spi_data_r[12] ;
    input \spi_data_r[13] ;
    input \spi_data_r[14] ;
    input \spi_data_r[15] ;
    input \spi_data_r[16] ;
    input \spi_data_r[17] ;
    input \spi_data_r[18] ;
    input \spi_data_r[19] ;
    input \spi_data_r[20] ;
    input \spi_data_r[21] ;
    input \spi_data_r[22] ;
    input \spi_data_r[23] ;
    input \spi_data_r[24] ;
    input \spi_data_r[25] ;
    input \spi_data_r[26] ;
    input \spi_data_r[27] ;
    input \spi_data_r[28] ;
    input \spi_data_r[29] ;
    input \spi_data_r[30] ;
    input \spi_data_r[31] ;
    output \quad_homing[1] ;
    input clk_enable_505;
    input n29120;
    input n13052;
    input n26969;
    input pin_io_out_34;
    output n27632;
    
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire [1:0]sync /* synthesis ASYNC_REG="TRUE" */ ;   // c:/s_links/sources/quad_decoder.v(106[30:34])
    wire [1:0]AB /* synthesis ASYNC_REG="TRUE" */ ;   // c:/s_links/sources/quad_decoder.v(106[36:38])
    wire \pin_intrpt[11]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[11] */ ;   // c:/s_links/sources/mcm_top.v(102[46:56])
    
    wire clk_1MHz_enable_246, n26155;
    wire [31:0]quad_set;   // c:/s_links/sources/quad_decoder.v(40[31:39])
    wire [1:0]quad_homing;   // c:/s_links/sources/quad_decoder.v(41[19:30])
    wire [3:0]n1901;
    
    wire n28793, n9639, n26749, n9647, n9652, quad_set_valid, spi_data_out_r_39__N_1864, 
        n10928, n25190, n11542;
    wire [31:0]n6236;
    
    wire n25189, n25188, n25187, n25186, n25185, n25184, n25183, 
        n25182, n25181, n25180, n25179, n25178, n25177, n3, n27025, 
        n25833, n25831, n25853, n25851, n25176, n25873, n25871, 
        n25893, n25175, n25891, n25913, n25911, n25933, n25931, 
        n25953, n25951, n25973, n25971, n25993, n25991, n26013, 
        n26011, n26033, n26031, n26061, n26059, n26087, n26085, 
        n26107, n26105, n26135, n26133, n26165, n28717, n28716, 
        n4, n27;
    
    FD1P3AX quad_count_i0_i0 (.D(n26155), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_1781[0] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX sync_i0 (.D(\quad_b[3] ), .CK(clk_1MHz), .Q(sync[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam sync_i0.GSR = "DISABLED";
    FD1S3AX AB_i0 (.D(sync[0]), .CK(clk_1MHz), .Q(AB[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam AB_i0.GSR = "DISABLED";
    FD1S3AX quad_buffer_i0 (.D(quad_count[0]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i0.GSR = "DISABLED";
    FD1P3IX quad_set__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i0.GSR = "DISABLED";
    FD1P3IX quad_homing__i0 (.D(n29762), .SP(clk_enable_434), .CD(n29239), 
            .CK(clk), .Q(quad_homing[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam quad_homing__i0.GSR = "DISABLED";
    FD1S3JX state_FSM_i0 (.D(n28793), .CK(clk_1MHz), .PD(n29239), .Q(n1901[0]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i0.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut (.A(n1901[3]), .B(AB[1]), .C(AB[0]), .D(n9639), 
         .Z(n26749)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i1_4_lut_4_lut.init = 16'h96c3;
    LUT4 i4868_4_lut_4_lut (.A(n1901[2]), .B(AB[0]), .C(AB[1]), .D(n9647), 
         .Z(n9652)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C (D))))) */ ;   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam i4868_4_lut_4_lut.init = 16'h3828;
    FD1S3IX quad_set_complete_451 (.D(quad_set_valid), .CK(clk_1MHz), .CD(n29239), 
            .Q(quad_set_complete)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_set_complete_451.GSR = "DISABLED";
    FD1S3IX i41_407 (.D(spi_data_out_r_39__N_1864), .CK(clk), .CD(n29239), 
            .Q(spi_data_out_r_39__N_1676)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam i41_407.GSR = "DISABLED";
    LUT4 i4678_4_lut (.A(AB[0]), .B(AB[1]), .C(n1901[2]), .D(n1901[1]), 
         .Z(n10928)) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A (B+!(C))) */ ;
    defparam i4678_4_lut.init = 16'he7ed;
    LUT4 i22607_2_lut_2_lut_4_lut (.A(n29098), .B(\spi_addr[0] ), .C(n26933), 
         .D(n13511), .Z(spi_data_out_r_39__N_2332)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (D))) */ ;
    defparam i22607_2_lut_2_lut_4_lut.init = 16'h005d;
    LUT4 i22592_2_lut_2_lut_4_lut (.A(n29098), .B(\spi_addr[0] ), .C(n26933), 
         .D(n13506), .Z(spi_data_out_r_39__N_1396)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (D))) */ ;
    defparam i22592_2_lut_2_lut_4_lut.init = 16'h005d;
    LUT4 i22598_2_lut_2_lut_4_lut (.A(n29098), .B(\spi_addr[0] ), .C(n26933), 
         .D(n13413), .Z(spi_data_out_r_39__N_1864)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (D))) */ ;
    defparam i22598_2_lut_2_lut_4_lut.init = 16'h005d;
    FD1S3AX quad_buffer_i31 (.D(quad_count[31]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i31.GSR = "DISABLED";
    FD1S3AX quad_buffer_i30 (.D(quad_count[30]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i30.GSR = "DISABLED";
    FD1S3AX quad_buffer_i29 (.D(quad_count[29]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i29.GSR = "DISABLED";
    FD1S3AX quad_buffer_i28 (.D(quad_count[28]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i28.GSR = "DISABLED";
    FD1S3AX quad_buffer_i27 (.D(quad_count[27]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i27.GSR = "DISABLED";
    FD1S3AX quad_buffer_i26 (.D(quad_count[26]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i26.GSR = "DISABLED";
    FD1S3AX quad_buffer_i25 (.D(quad_count[25]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i25.GSR = "DISABLED";
    FD1S3AX quad_buffer_i24 (.D(quad_count[24]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i24.GSR = "DISABLED";
    FD1S3AX quad_buffer_i23 (.D(quad_count[23]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i23.GSR = "DISABLED";
    FD1S3AX quad_buffer_i22 (.D(quad_count[22]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i22.GSR = "DISABLED";
    FD1S3AX quad_buffer_i21 (.D(quad_count[21]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i21.GSR = "DISABLED";
    FD1S3AX quad_buffer_i20 (.D(quad_count[20]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i20.GSR = "DISABLED";
    FD1S3AX quad_buffer_i19 (.D(quad_count[19]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i19.GSR = "DISABLED";
    FD1S3AX quad_buffer_i18 (.D(quad_count[18]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i18.GSR = "DISABLED";
    FD1S3AX quad_buffer_i17 (.D(quad_count[17]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i17.GSR = "DISABLED";
    FD1S3AX quad_buffer_i16 (.D(quad_count[16]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i16.GSR = "DISABLED";
    FD1S3AX quad_buffer_i15 (.D(quad_count[15]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i15.GSR = "DISABLED";
    FD1S3AX quad_buffer_i14 (.D(quad_count[14]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i14.GSR = "DISABLED";
    FD1S3AX quad_buffer_i13 (.D(quad_count[13]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i13.GSR = "DISABLED";
    FD1S3AX quad_buffer_i12 (.D(quad_count[12]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i12.GSR = "DISABLED";
    FD1S3AX quad_buffer_i11 (.D(quad_count[11]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i11.GSR = "DISABLED";
    FD1S3AX quad_buffer_i10 (.D(quad_count[10]), .CK(\pin_intrpt[11] ), 
            .Q(quad_buffer[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i10.GSR = "DISABLED";
    FD1S3AX quad_buffer_i9 (.D(quad_count[9]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i9.GSR = "DISABLED";
    FD1S3AX quad_buffer_i8 (.D(quad_count[8]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i8.GSR = "DISABLED";
    FD1S3AX quad_buffer_i7 (.D(quad_count[7]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i7.GSR = "DISABLED";
    FD1S3AX quad_buffer_i6 (.D(quad_count[6]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i6.GSR = "DISABLED";
    FD1S3AX quad_buffer_i5 (.D(quad_count[5]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i5.GSR = "DISABLED";
    FD1S3AX quad_buffer_i4 (.D(quad_count[4]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i4.GSR = "DISABLED";
    FD1S3AX quad_buffer_i3 (.D(quad_count[3]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i3.GSR = "DISABLED";
    FD1S3AX quad_buffer_i2 (.D(quad_count[2]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i2.GSR = "DISABLED";
    FD1S3AX quad_buffer_i1 (.D(quad_count[1]), .CK(\pin_intrpt[11] ), .Q(quad_buffer[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i1.GSR = "DISABLED";
    FD1S3AX AB_i1 (.D(sync[1]), .CK(clk_1MHz), .Q(AB[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam AB_i1.GSR = "DISABLED";
    FD1S3AX sync_i1 (.D(\quad_a[3] ), .CK(clk_1MHz), .Q(sync[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam sync_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_1781[31] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    CCU2D add_2013_33 (.A0(resetn_c), .B0(n11542), .C0(quad_count[30]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[31]), 
          .D1(GND_net), .CIN(n25190), .S0(n6236[30]), .S1(n6236[31]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_33.INIT0 = 16'hd2d2;
    defparam add_2013_33.INIT1 = 16'hd2d2;
    defparam add_2013_33.INJECT1_0 = "NO";
    defparam add_2013_33.INJECT1_1 = "NO";
    CCU2D add_2013_31 (.A0(resetn_c), .B0(n11542), .C0(quad_count[28]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[29]), 
          .D1(GND_net), .CIN(n25189), .COUT(n25190), .S0(n6236[28]), 
          .S1(n6236[29]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_31.INIT0 = 16'hd2d2;
    defparam add_2013_31.INIT1 = 16'hd2d2;
    defparam add_2013_31.INJECT1_0 = "NO";
    defparam add_2013_31.INJECT1_1 = "NO";
    FD1S3AX spi_data_out_r_i31 (.D(\spi_data_out_r_39__N_1781[30] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i30 (.D(\spi_data_out_r_39__N_1781[29] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i29 (.D(\spi_data_out_r_39__N_1781[28] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i28 (.D(\spi_data_out_r_39__N_1781[27] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i27 (.D(\spi_data_out_r_39__N_1781[26] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i26 (.D(\spi_data_out_r_39__N_1781[25] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    CCU2D add_2013_29 (.A0(resetn_c), .B0(n11542), .C0(quad_count[26]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[27]), 
          .D1(GND_net), .CIN(n25188), .COUT(n25189), .S0(n6236[26]), 
          .S1(n6236[27]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_29.INIT0 = 16'hd2d2;
    defparam add_2013_29.INIT1 = 16'hd2d2;
    defparam add_2013_29.INJECT1_0 = "NO";
    defparam add_2013_29.INJECT1_1 = "NO";
    CCU2D add_2013_27 (.A0(resetn_c), .B0(n11542), .C0(quad_count[24]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[25]), 
          .D1(GND_net), .CIN(n25187), .COUT(n25188), .S0(n6236[24]), 
          .S1(n6236[25]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_27.INIT0 = 16'hd2d2;
    defparam add_2013_27.INIT1 = 16'hd2d2;
    defparam add_2013_27.INJECT1_0 = "NO";
    defparam add_2013_27.INJECT1_1 = "NO";
    CCU2D add_2013_25 (.A0(resetn_c), .B0(n11542), .C0(quad_count[22]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[23]), 
          .D1(GND_net), .CIN(n25186), .COUT(n25187), .S0(n6236[22]), 
          .S1(n6236[23]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_25.INIT0 = 16'hd2d2;
    defparam add_2013_25.INIT1 = 16'hd2d2;
    defparam add_2013_25.INJECT1_0 = "NO";
    defparam add_2013_25.INJECT1_1 = "NO";
    CCU2D add_2013_23 (.A0(resetn_c), .B0(n11542), .C0(quad_count[20]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[21]), 
          .D1(GND_net), .CIN(n25185), .COUT(n25186), .S0(n6236[20]), 
          .S1(n6236[21]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_23.INIT0 = 16'hd2d2;
    defparam add_2013_23.INIT1 = 16'hd2d2;
    defparam add_2013_23.INJECT1_0 = "NO";
    defparam add_2013_23.INJECT1_1 = "NO";
    CCU2D add_2013_21 (.A0(resetn_c), .B0(n11542), .C0(quad_count[18]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[19]), 
          .D1(GND_net), .CIN(n25184), .COUT(n25185), .S0(n6236[18]), 
          .S1(n6236[19]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_21.INIT0 = 16'hd2d2;
    defparam add_2013_21.INIT1 = 16'hd2d2;
    defparam add_2013_21.INJECT1_0 = "NO";
    defparam add_2013_21.INJECT1_1 = "NO";
    CCU2D add_2013_19 (.A0(resetn_c), .B0(n11542), .C0(quad_count[16]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[17]), 
          .D1(GND_net), .CIN(n25183), .COUT(n25184), .S0(n6236[16]), 
          .S1(n6236[17]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_19.INIT0 = 16'hd2d2;
    defparam add_2013_19.INIT1 = 16'hd2d2;
    defparam add_2013_19.INJECT1_0 = "NO";
    defparam add_2013_19.INJECT1_1 = "NO";
    FD1S3AX spi_data_out_r_i25 (.D(\spi_data_out_r_39__N_1781[24] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i24 (.D(\spi_data_out_r_39__N_1781[23] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i23 (.D(\spi_data_out_r_39__N_1781[22] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i22 (.D(\spi_data_out_r_39__N_1781[21] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i21 (.D(\spi_data_out_r_39__N_1781[20] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i20 (.D(\spi_data_out_r_39__N_1781[19] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i19 (.D(\spi_data_out_r_39__N_1781[18] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i18 (.D(\spi_data_out_r_39__N_1781[17] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i17 (.D(\spi_data_out_r_39__N_1781[16] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i16 (.D(\spi_data_out_r_39__N_1781[15] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_1781[14] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_1781[13] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_1781[12] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_1781[11] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_1781[10] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_1781[9] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_1781[8] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_1781[7] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_1781[6] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_1781[5] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_1781[4] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    CCU2D add_2013_17 (.A0(resetn_c), .B0(n11542), .C0(quad_count[14]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[15]), 
          .D1(GND_net), .CIN(n25182), .COUT(n25183), .S0(n6236[14]), 
          .S1(n6236[15]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_17.INIT0 = 16'hd2d2;
    defparam add_2013_17.INIT1 = 16'hd2d2;
    defparam add_2013_17.INJECT1_0 = "NO";
    defparam add_2013_17.INJECT1_1 = "NO";
    CCU2D add_2013_15 (.A0(resetn_c), .B0(n11542), .C0(quad_count[12]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[13]), 
          .D1(GND_net), .CIN(n25181), .COUT(n25182), .S0(n6236[12]), 
          .S1(n6236[13]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_15.INIT0 = 16'hd2d2;
    defparam add_2013_15.INIT1 = 16'hd2d2;
    defparam add_2013_15.INJECT1_0 = "NO";
    defparam add_2013_15.INJECT1_1 = "NO";
    CCU2D add_2013_13 (.A0(resetn_c), .B0(n11542), .C0(quad_count[10]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[11]), 
          .D1(GND_net), .CIN(n25180), .COUT(n25181), .S0(n6236[10]), 
          .S1(n6236[11]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_13.INIT0 = 16'hd2d2;
    defparam add_2013_13.INIT1 = 16'hd2d2;
    defparam add_2013_13.INJECT1_0 = "NO";
    defparam add_2013_13.INJECT1_1 = "NO";
    CCU2D add_2013_11 (.A0(resetn_c), .B0(n11542), .C0(quad_count[8]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[9]), 
          .D1(GND_net), .CIN(n25179), .COUT(n25180), .S0(n6236[8]), 
          .S1(n6236[9]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_11.INIT0 = 16'hd2d2;
    defparam add_2013_11.INIT1 = 16'hd2d2;
    defparam add_2013_11.INJECT1_0 = "NO";
    defparam add_2013_11.INJECT1_1 = "NO";
    CCU2D add_2013_9 (.A0(resetn_c), .B0(n11542), .C0(quad_count[6]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[7]), 
          .D1(GND_net), .CIN(n25178), .COUT(n25179), .S0(n6236[6]), 
          .S1(n6236[7]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_9.INIT0 = 16'hd2d2;
    defparam add_2013_9.INIT1 = 16'hd2d2;
    defparam add_2013_9.INJECT1_0 = "NO";
    defparam add_2013_9.INJECT1_1 = "NO";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_1781[3] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_1781[2] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_1781[1] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1636[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    CCU2D add_2013_7 (.A0(resetn_c), .B0(n11542), .C0(quad_count[4]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[5]), 
          .D1(GND_net), .CIN(n25177), .COUT(n25178), .S0(n6236[4]), 
          .S1(n6236[5]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_7.INIT0 = 16'hd2d2;
    defparam add_2013_7.INIT1 = 16'hd2d2;
    defparam add_2013_7.INJECT1_0 = "NO";
    defparam add_2013_7.INJECT1_1 = "NO";
    LUT4 i31_4_lut (.A(n6236[31]), .B(quad_set[31]), .C(n3), .D(n27025), 
         .Z(n25833)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut.init = 16'hcac0;
    LUT4 i31_4_lut_adj_871 (.A(n6236[30]), .B(quad_set[30]), .C(n3), .D(n27025), 
         .Z(n25831)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_871.init = 16'hcac0;
    LUT4 i31_4_lut_adj_872 (.A(n6236[29]), .B(quad_set[29]), .C(n3), .D(n27025), 
         .Z(n25853)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_872.init = 16'hcac0;
    LUT4 i31_4_lut_adj_873 (.A(n6236[28]), .B(quad_set[28]), .C(n3), .D(n27025), 
         .Z(n25851)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_873.init = 16'hcac0;
    CCU2D add_2013_5 (.A0(resetn_c), .B0(n11542), .C0(quad_count[2]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[3]), 
          .D1(GND_net), .CIN(n25176), .COUT(n25177), .S0(n6236[2]), 
          .S1(n6236[3]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_5.INIT0 = 16'hd2d2;
    defparam add_2013_5.INIT1 = 16'hd2d2;
    defparam add_2013_5.INJECT1_0 = "NO";
    defparam add_2013_5.INJECT1_1 = "NO";
    LUT4 i31_4_lut_adj_874 (.A(n6236[27]), .B(quad_set[27]), .C(n3), .D(n27025), 
         .Z(n25873)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_874.init = 16'hcac0;
    LUT4 i31_4_lut_adj_875 (.A(n6236[26]), .B(quad_set[26]), .C(n3), .D(n27025), 
         .Z(n25871)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_875.init = 16'hcac0;
    LUT4 i31_4_lut_adj_876 (.A(n6236[25]), .B(quad_set[25]), .C(n3), .D(n27025), 
         .Z(n25893)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_876.init = 16'hcac0;
    CCU2D add_2013_3 (.A0(resetn_c), .B0(n11542), .C0(quad_count[0]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11542), .C1(quad_count[1]), 
          .D1(GND_net), .CIN(n25175), .COUT(n25176), .S0(n6236[0]), 
          .S1(n6236[1]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_3.INIT0 = 16'h2d2d;
    defparam add_2013_3.INIT1 = 16'hd2d2;
    defparam add_2013_3.INJECT1_0 = "NO";
    defparam add_2013_3.INJECT1_1 = "NO";
    LUT4 i31_4_lut_adj_877 (.A(n6236[24]), .B(quad_set[24]), .C(n3), .D(n27025), 
         .Z(n25891)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_877.init = 16'hcac0;
    LUT4 i31_4_lut_adj_878 (.A(n6236[23]), .B(quad_set[23]), .C(n3), .D(n27025), 
         .Z(n25913)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_878.init = 16'hcac0;
    FD1P3AX quad_count_i0_i31 (.D(n25833), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i31.GSR = "DISABLED";
    LUT4 i31_4_lut_adj_879 (.A(n6236[22]), .B(quad_set[22]), .C(n3), .D(n27025), 
         .Z(n25911)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_879.init = 16'hcac0;
    FD1P3AX quad_count_i0_i30 (.D(n25831), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i30.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i29 (.D(n25853), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i29.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i28 (.D(n25851), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i28.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i27 (.D(n25873), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i27.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i26 (.D(n25871), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i26.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i25 (.D(n25893), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i25.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i24 (.D(n25891), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i24.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i23 (.D(n25913), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i23.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i22 (.D(n25911), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i22.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i21 (.D(n25933), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i21.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i20 (.D(n25931), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i20.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i19 (.D(n25953), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i19.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i18 (.D(n25951), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i18.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i17 (.D(n25973), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i17.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i16 (.D(n25971), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i16.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i15 (.D(n25993), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i15.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i14 (.D(n25991), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i14.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i13 (.D(n26013), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i13.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i12 (.D(n26011), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i12.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i11 (.D(n26033), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i11.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i10 (.D(n26031), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i10.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i9 (.D(n26061), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i9.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i8 (.D(n26059), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i8.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i7 (.D(n26087), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i7.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i6 (.D(n26085), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i6.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i5 (.D(n26107), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i5.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i4 (.D(n26105), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i4.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i3 (.D(n26135), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i3.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i2 (.D(n26133), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i1 (.D(n26165), .SP(clk_1MHz_enable_246), .CK(clk_1MHz), 
            .Q(quad_count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i1.GSR = "DISABLED";
    LUT4 i31_4_lut_adj_880 (.A(n6236[21]), .B(quad_set[21]), .C(n3), .D(n27025), 
         .Z(n25933)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_880.init = 16'hcac0;
    LUT4 i4679_3_lut_4_lut (.A(AB[0]), .B(AB[1]), .C(n1901[3]), .D(n10928), 
         .Z(n11542)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // c:/s_links/sources/quad_decoder.v(162[19:30])
    defparam i4679_3_lut_4_lut.init = 16'hbfb0;
    CCU2D add_2013_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(resetn_c), .B1(n11542), .C1(GND_net), .D1(GND_net), .COUT(n25175));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2013_1.INIT0 = 16'hF000;
    defparam add_2013_1.INIT1 = 16'hdddd;
    defparam add_2013_1.INJECT1_0 = "NO";
    defparam add_2013_1.INJECT1_1 = "NO";
    LUT4 i31_4_lut_adj_881 (.A(n6236[20]), .B(quad_set[20]), .C(n3), .D(n27025), 
         .Z(n25931)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_881.init = 16'hcac0;
    LUT4 i31_4_lut_adj_882 (.A(n6236[19]), .B(quad_set[19]), .C(n3), .D(n27025), 
         .Z(n25953)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_882.init = 16'hcac0;
    LUT4 i31_4_lut_adj_883 (.A(n6236[18]), .B(quad_set[18]), .C(n3), .D(n27025), 
         .Z(n25951)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_883.init = 16'hcac0;
    LUT4 i31_4_lut_adj_884 (.A(n6236[17]), .B(quad_set[17]), .C(n3), .D(n27025), 
         .Z(n25973)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_884.init = 16'hcac0;
    LUT4 i31_4_lut_adj_885 (.A(n6236[16]), .B(quad_set[16]), .C(n3), .D(n27025), 
         .Z(n25971)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_885.init = 16'hcac0;
    LUT4 i31_4_lut_adj_886 (.A(n6236[15]), .B(quad_set[15]), .C(n3), .D(n27025), 
         .Z(n25993)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_886.init = 16'hcac0;
    LUT4 i31_4_lut_adj_887 (.A(n6236[14]), .B(quad_set[14]), .C(n3), .D(n27025), 
         .Z(n25991)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_887.init = 16'hcac0;
    LUT4 i31_4_lut_adj_888 (.A(n6236[13]), .B(quad_set[13]), .C(n3), .D(n27025), 
         .Z(n26013)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_888.init = 16'hcac0;
    LUT4 i31_4_lut_adj_889 (.A(n6236[12]), .B(quad_set[12]), .C(n3), .D(n27025), 
         .Z(n26011)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_889.init = 16'hcac0;
    LUT4 i31_4_lut_adj_890 (.A(n6236[11]), .B(quad_set[11]), .C(n3), .D(n27025), 
         .Z(n26033)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_890.init = 16'hcac0;
    LUT4 i31_4_lut_adj_891 (.A(n6236[10]), .B(quad_set[10]), .C(n3), .D(n27025), 
         .Z(n26031)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_891.init = 16'hcac0;
    LUT4 i31_4_lut_adj_892 (.A(n6236[9]), .B(quad_set[9]), .C(n3), .D(n27025), 
         .Z(n26061)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_892.init = 16'hcac0;
    LUT4 i31_4_lut_adj_893 (.A(n6236[8]), .B(quad_set[8]), .C(n3), .D(n27025), 
         .Z(n26059)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_893.init = 16'hcac0;
    LUT4 i31_4_lut_adj_894 (.A(n6236[7]), .B(quad_set[7]), .C(n3), .D(n27025), 
         .Z(n26087)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_894.init = 16'hcac0;
    LUT4 i31_4_lut_adj_895 (.A(n6236[6]), .B(quad_set[6]), .C(n3), .D(n27025), 
         .Z(n26085)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_895.init = 16'hcac0;
    LUT4 i31_4_lut_adj_896 (.A(n6236[5]), .B(quad_set[5]), .C(n3), .D(n27025), 
         .Z(n26107)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_896.init = 16'hcac0;
    LUT4 i31_4_lut_adj_897 (.A(n6236[4]), .B(quad_set[4]), .C(n3), .D(n27025), 
         .Z(n26105)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_897.init = 16'hcac0;
    LUT4 i31_4_lut_adj_898 (.A(n6236[3]), .B(quad_set[3]), .C(n3), .D(n27025), 
         .Z(n26135)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_898.init = 16'hcac0;
    LUT4 i31_4_lut_adj_899 (.A(n6236[2]), .B(quad_set[2]), .C(n3), .D(n27025), 
         .Z(n26133)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_899.init = 16'hcac0;
    LUT4 i31_4_lut_adj_900 (.A(n6236[1]), .B(quad_set[1]), .C(n3), .D(n27025), 
         .Z(n26165)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_900.init = 16'hcac0;
    FD1P3IX quad_set__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i1.GSR = "DISABLED";
    FD1P3IX quad_set__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i2.GSR = "DISABLED";
    FD1P3IX quad_set__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i3.GSR = "DISABLED";
    FD1P3IX quad_set__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i4.GSR = "DISABLED";
    FD1P3IX quad_set__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i5.GSR = "DISABLED";
    FD1P3IX quad_set__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i6.GSR = "DISABLED";
    FD1P3IX quad_set__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i7.GSR = "DISABLED";
    FD1P3IX quad_set__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i8.GSR = "DISABLED";
    FD1P3IX quad_set__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i9.GSR = "DISABLED";
    FD1P3IX quad_set__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i10.GSR = "DISABLED";
    FD1P3IX quad_set__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i11.GSR = "DISABLED";
    FD1P3IX quad_set__i12 (.D(\spi_data_r[12] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i12.GSR = "DISABLED";
    FD1P3IX quad_set__i13 (.D(\spi_data_r[13] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i13.GSR = "DISABLED";
    FD1P3IX quad_set__i14 (.D(\spi_data_r[14] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i14.GSR = "DISABLED";
    FD1P3IX quad_set__i15 (.D(\spi_data_r[15] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i15.GSR = "DISABLED";
    FD1P3IX quad_set__i16 (.D(\spi_data_r[16] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i16.GSR = "DISABLED";
    FD1P3IX quad_set__i17 (.D(\spi_data_r[17] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i17.GSR = "DISABLED";
    FD1P3IX quad_set__i18 (.D(\spi_data_r[18] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i18.GSR = "DISABLED";
    FD1P3IX quad_set__i19 (.D(\spi_data_r[19] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i19.GSR = "DISABLED";
    FD1P3IX quad_set__i20 (.D(\spi_data_r[20] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i20.GSR = "DISABLED";
    FD1P3IX quad_set__i21 (.D(\spi_data_r[21] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i21.GSR = "DISABLED";
    FD1P3IX quad_set__i22 (.D(\spi_data_r[22] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i22.GSR = "DISABLED";
    FD1P3IX quad_set__i23 (.D(\spi_data_r[23] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i23.GSR = "DISABLED";
    FD1P3IX quad_set__i24 (.D(\spi_data_r[24] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i24.GSR = "DISABLED";
    FD1P3IX quad_set__i25 (.D(\spi_data_r[25] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i25.GSR = "DISABLED";
    FD1P3IX quad_set__i26 (.D(\spi_data_r[26] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i26.GSR = "DISABLED";
    FD1P3IX quad_set__i27 (.D(\spi_data_r[27] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i27.GSR = "DISABLED";
    FD1P3IX quad_set__i28 (.D(\spi_data_r[28] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i28.GSR = "DISABLED";
    FD1P3IX quad_set__i29 (.D(\spi_data_r[29] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i29.GSR = "DISABLED";
    FD1P3IX quad_set__i30 (.D(\spi_data_r[30] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i30.GSR = "DISABLED";
    FD1P3IX quad_set__i31 (.D(\spi_data_r[31] ), .SP(clk_enable_398), .CD(n29239), 
            .CK(clk), .Q(quad_set[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i31.GSR = "DISABLED";
    FD1P3IX quad_homing__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_434), .CD(n29239), 
            .CK(clk), .Q(\quad_homing[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam quad_homing__i1.GSR = "DISABLED";
    FD1S3IX state_FSM_i1 (.D(n28717), .CK(clk_1MHz), .CD(n29239), .Q(n1901[1]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i1.GSR = "DISABLED";
    FD1S3IX state_FSM_i2 (.D(n9652), .CK(clk_1MHz), .CD(n29239), .Q(n1901[2]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i2.GSR = "DISABLED";
    FD1S3IX state_FSM_i3 (.D(n28716), .CK(clk_1MHz), .CD(n29239), .Q(n1901[3]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i3.GSR = "DISABLED";
    FD1P3IX quad_set_valid_404 (.D(n29120), .SP(clk_enable_505), .CD(n29239), 
            .CK(clk), .Q(quad_set_valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set_valid_404.GSR = "DISABLED";
    LUT4 AB_1__bdd_4_lut_23071 (.A(AB[1]), .B(n1901[1]), .C(AB[0]), .D(n9647), 
         .Z(n28717)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B (C (D))))) */ ;
    defparam AB_1__bdd_4_lut_23071.init = 16'h5848;
    LUT4 AB_1__bdd_4_lut_23035 (.A(AB[1]), .B(n1901[3]), .C(AB[0]), .D(n9639), 
         .Z(n28716)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam AB_1__bdd_4_lut_23035.init = 16'ha484;
    LUT4 AB_1__bdd_4_lut (.A(AB[1]), .B(n1901[0]), .C(AB[0]), .D(n9639), 
         .Z(n28793)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B (C+!(D)))) */ ;
    defparam AB_1__bdd_4_lut.init = 16'h8584;
    LUT4 reduce_or_501_i1_2_lut (.A(n1901[3]), .B(n1901[0]), .Z(n9647)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam reduce_or_501_i1_2_lut.init = 16'heeee;
    LUT4 i22912_4_lut (.A(quad_set_valid), .B(resetn_c), .C(n26749), .D(n13052), 
         .Z(clk_1MHz_enable_246)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i22912_4_lut.init = 16'hffbf;
    LUT4 i31_4_lut_adj_901 (.A(n6236[0]), .B(quad_set[0]), .C(n3), .D(n27025), 
         .Z(n26155)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_901.init = 16'hcac0;
    LUT4 i3_4_lut (.A(quad_set_valid), .B(n26969), .C(resetn_c), .D(n4), 
         .Z(n3)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i1_3_lut (.A(resetn_c), .B(n13052), .C(n4), .Z(n27025)) /* synthesis lut_function=(!((B (C))+!A)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i1_3_lut.init = 16'h2a2a;
    LUT4 i1_4_lut (.A(n1901[1]), .B(n27), .C(n1901[2]), .D(n1901[3]), 
         .Z(n4)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i1_4_lut.init = 16'h33c9;
    LUT4 i15_2_lut (.A(AB[1]), .B(AB[0]), .Z(n27)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(155[16] 158[10])
    defparam i15_2_lut.init = 16'h6666;
    LUT4 i22462_2_lut (.A(quad_homing[0]), .B(pin_io_out_34), .Z(n27632)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22462_2_lut.init = 16'h8888;
    LUT4 reduce_or_506_i1_2_lut (.A(n1901[2]), .B(n1901[1]), .Z(n9639)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam reduce_or_506_i1_2_lut.init = 16'heeee;
    
endmodule
//
// Verilog Description of module \servo(DEV_ID=6,UART_ADDRESS_WIDTH=4) 
//

module \servo(DEV_ID=6,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_170, 
            n29239, \spi_data_r[0] , n29191, n29196, mode_adj_182, 
            n14, C_5_c_c, n29267, n8633) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_170;
    input n29239;
    input \spi_data_r[0] ;
    input n29191;
    input n29196;
    input mode_adj_182;
    output n14;
    input C_5_c_c;
    input n29267;
    output n8633;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    FD1P3IX mode_60 (.D(\spi_data_r[0] ), .SP(clk_enable_170), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=418, LSE_RLINE=453 */ ;   // c:/s_links/sources/slot_cards/servo.v(66[8] 74[4])
    defparam mode_60.GSR = "DISABLED";
    LUT4 i2_2_lut_3_lut_4_lut (.A(mode), .B(n29191), .C(n29196), .D(mode_adj_182), 
         .Z(n14)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (C+!(D)))) */ ;   // c:/s_links/sources/slot_cards/servo.v(61[19:72])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h2f22;
    LUT4 i22845_3_lut_4_lut (.A(mode), .B(n29191), .C(C_5_c_c), .D(n29267), 
         .Z(n8633)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;   // c:/s_links/sources/slot_cards/servo.v(61[19:72])
    defparam i22845_3_lut_4_lut.init = 16'hfd00;
    
endmodule
//
// Verilog Description of module \quad_decoder(DEV_ID=4) 
//

module \quad_decoder(DEV_ID=4)  (quad_count, clk_1MHz, \spi_data_out_r_39__N_1870[0] , 
            clk, \spi_data_out_r_39__N_2015[0] , \quad_b[4] , quad_buffer, 
            \pin_intrpt[14] , n29239, clk_enable_162, \spi_data_r[0] , 
            quad_homing, clk_enable_77, n29762, \spi_data_r[1] , \spi_data_r[31] , 
            \spi_data_r[30] , \spi_data_r[29] , \spi_data_r[28] , \spi_data_r[27] , 
            \spi_data_r[26] , \spi_data_r[25] , \spi_data_r[24] , \spi_data_r[23] , 
            \spi_data_r[22] , \spi_data_r[21] , \spi_data_r[20] , \spi_data_r[19] , 
            \spi_data_r[18] , \spi_data_r[17] , \spi_data_r[16] , \spi_data_r[15] , 
            \spi_data_r[14] , \spi_data_r[13] , \spi_data_r[12] , \spi_data_r[11] , 
            \spi_data_r[10] , \spi_data_r[9] , \spi_data_r[8] , \spi_data_r[7] , 
            \spi_data_r[6] , \spi_data_r[5] , \spi_data_r[4] , \spi_data_r[3] , 
            \spi_data_r[2] , quad_set_complete, spi_data_out_r_39__N_1910, 
            spi_data_out_r_39__N_2098, \quad_a[4] , \spi_data_out_r_39__N_1870[31] , 
            \spi_data_out_r_39__N_2015[31] , \spi_data_out_r_39__N_1870[30] , 
            \spi_data_out_r_39__N_2015[30] , \spi_data_out_r_39__N_1870[29] , 
            \spi_data_out_r_39__N_2015[29] , \spi_data_out_r_39__N_1870[28] , 
            \spi_data_out_r_39__N_2015[28] , \spi_data_out_r_39__N_1870[27] , 
            \spi_data_out_r_39__N_2015[27] , \spi_data_out_r_39__N_1870[26] , 
            \spi_data_out_r_39__N_2015[26] , \spi_data_out_r_39__N_1870[25] , 
            \spi_data_out_r_39__N_2015[25] , \spi_data_out_r_39__N_1870[24] , 
            \spi_data_out_r_39__N_2015[24] , \spi_data_out_r_39__N_1870[23] , 
            \spi_data_out_r_39__N_2015[23] , \spi_data_out_r_39__N_1870[22] , 
            \spi_data_out_r_39__N_2015[22] , \spi_data_out_r_39__N_1870[21] , 
            \spi_data_out_r_39__N_2015[21] , \spi_data_out_r_39__N_1870[20] , 
            \spi_data_out_r_39__N_2015[20] , \spi_data_out_r_39__N_1870[19] , 
            \spi_data_out_r_39__N_2015[19] , \spi_data_out_r_39__N_1870[18] , 
            \spi_data_out_r_39__N_2015[18] , \spi_data_out_r_39__N_1870[17] , 
            \spi_data_out_r_39__N_2015[17] , \spi_data_out_r_39__N_1870[16] , 
            \spi_data_out_r_39__N_2015[16] , \spi_data_out_r_39__N_1870[15] , 
            \spi_data_out_r_39__N_2015[15] , \spi_data_out_r_39__N_1870[14] , 
            \spi_data_out_r_39__N_2015[14] , \spi_data_out_r_39__N_1870[13] , 
            \spi_data_out_r_39__N_2015[13] , \spi_data_out_r_39__N_1870[12] , 
            \spi_data_out_r_39__N_2015[12] , \spi_data_out_r_39__N_1870[11] , 
            \spi_data_out_r_39__N_2015[11] , \spi_data_out_r_39__N_1870[10] , 
            \spi_data_out_r_39__N_2015[10] , \spi_data_out_r_39__N_1870[9] , 
            \spi_data_out_r_39__N_2015[9] , \spi_data_out_r_39__N_1870[8] , 
            \spi_data_out_r_39__N_2015[8] , \spi_data_out_r_39__N_1870[7] , 
            \spi_data_out_r_39__N_2015[7] , \spi_data_out_r_39__N_1870[6] , 
            \spi_data_out_r_39__N_2015[6] , \spi_data_out_r_39__N_1870[5] , 
            \spi_data_out_r_39__N_2015[5] , \spi_data_out_r_39__N_1870[4] , 
            \spi_data_out_r_39__N_2015[4] , \spi_data_out_r_39__N_1870[3] , 
            \spi_data_out_r_39__N_2015[3] , \spi_data_out_r_39__N_1870[2] , 
            \spi_data_out_r_39__N_2015[2] , \spi_data_out_r_39__N_1870[1] , 
            \spi_data_out_r_39__N_2015[1] , resetn_c, GND_net, clk_enable_518, 
            n29080, n26938) /* synthesis syn_module_defined=1 */ ;
    output [31:0]quad_count;
    input clk_1MHz;
    output \spi_data_out_r_39__N_1870[0] ;
    input clk;
    input \spi_data_out_r_39__N_2015[0] ;
    input \quad_b[4] ;
    output [31:0]quad_buffer;
    input \pin_intrpt[14] ;
    input n29239;
    input clk_enable_162;
    input \spi_data_r[0] ;
    output [1:0]quad_homing;
    input clk_enable_77;
    input n29762;
    input \spi_data_r[1] ;
    input \spi_data_r[31] ;
    input \spi_data_r[30] ;
    input \spi_data_r[29] ;
    input \spi_data_r[28] ;
    input \spi_data_r[27] ;
    input \spi_data_r[26] ;
    input \spi_data_r[25] ;
    input \spi_data_r[24] ;
    input \spi_data_r[23] ;
    input \spi_data_r[22] ;
    input \spi_data_r[21] ;
    input \spi_data_r[20] ;
    input \spi_data_r[19] ;
    input \spi_data_r[18] ;
    input \spi_data_r[17] ;
    input \spi_data_r[16] ;
    input \spi_data_r[15] ;
    input \spi_data_r[14] ;
    input \spi_data_r[13] ;
    input \spi_data_r[12] ;
    input \spi_data_r[11] ;
    input \spi_data_r[10] ;
    input \spi_data_r[9] ;
    input \spi_data_r[8] ;
    input \spi_data_r[7] ;
    input \spi_data_r[6] ;
    input \spi_data_r[5] ;
    input \spi_data_r[4] ;
    input \spi_data_r[3] ;
    input \spi_data_r[2] ;
    output quad_set_complete;
    output spi_data_out_r_39__N_1910;
    input spi_data_out_r_39__N_2098;
    input \quad_a[4] ;
    output \spi_data_out_r_39__N_1870[31] ;
    input \spi_data_out_r_39__N_2015[31] ;
    output \spi_data_out_r_39__N_1870[30] ;
    input \spi_data_out_r_39__N_2015[30] ;
    output \spi_data_out_r_39__N_1870[29] ;
    input \spi_data_out_r_39__N_2015[29] ;
    output \spi_data_out_r_39__N_1870[28] ;
    input \spi_data_out_r_39__N_2015[28] ;
    output \spi_data_out_r_39__N_1870[27] ;
    input \spi_data_out_r_39__N_2015[27] ;
    output \spi_data_out_r_39__N_1870[26] ;
    input \spi_data_out_r_39__N_2015[26] ;
    output \spi_data_out_r_39__N_1870[25] ;
    input \spi_data_out_r_39__N_2015[25] ;
    output \spi_data_out_r_39__N_1870[24] ;
    input \spi_data_out_r_39__N_2015[24] ;
    output \spi_data_out_r_39__N_1870[23] ;
    input \spi_data_out_r_39__N_2015[23] ;
    output \spi_data_out_r_39__N_1870[22] ;
    input \spi_data_out_r_39__N_2015[22] ;
    output \spi_data_out_r_39__N_1870[21] ;
    input \spi_data_out_r_39__N_2015[21] ;
    output \spi_data_out_r_39__N_1870[20] ;
    input \spi_data_out_r_39__N_2015[20] ;
    output \spi_data_out_r_39__N_1870[19] ;
    input \spi_data_out_r_39__N_2015[19] ;
    output \spi_data_out_r_39__N_1870[18] ;
    input \spi_data_out_r_39__N_2015[18] ;
    output \spi_data_out_r_39__N_1870[17] ;
    input \spi_data_out_r_39__N_2015[17] ;
    output \spi_data_out_r_39__N_1870[16] ;
    input \spi_data_out_r_39__N_2015[16] ;
    output \spi_data_out_r_39__N_1870[15] ;
    input \spi_data_out_r_39__N_2015[15] ;
    output \spi_data_out_r_39__N_1870[14] ;
    input \spi_data_out_r_39__N_2015[14] ;
    output \spi_data_out_r_39__N_1870[13] ;
    input \spi_data_out_r_39__N_2015[13] ;
    output \spi_data_out_r_39__N_1870[12] ;
    input \spi_data_out_r_39__N_2015[12] ;
    output \spi_data_out_r_39__N_1870[11] ;
    input \spi_data_out_r_39__N_2015[11] ;
    output \spi_data_out_r_39__N_1870[10] ;
    input \spi_data_out_r_39__N_2015[10] ;
    output \spi_data_out_r_39__N_1870[9] ;
    input \spi_data_out_r_39__N_2015[9] ;
    output \spi_data_out_r_39__N_1870[8] ;
    input \spi_data_out_r_39__N_2015[8] ;
    output \spi_data_out_r_39__N_1870[7] ;
    input \spi_data_out_r_39__N_2015[7] ;
    output \spi_data_out_r_39__N_1870[6] ;
    input \spi_data_out_r_39__N_2015[6] ;
    output \spi_data_out_r_39__N_1870[5] ;
    input \spi_data_out_r_39__N_2015[5] ;
    output \spi_data_out_r_39__N_1870[4] ;
    input \spi_data_out_r_39__N_2015[4] ;
    output \spi_data_out_r_39__N_1870[3] ;
    input \spi_data_out_r_39__N_2015[3] ;
    output \spi_data_out_r_39__N_1870[2] ;
    input \spi_data_out_r_39__N_2015[2] ;
    output \spi_data_out_r_39__N_1870[1] ;
    input \spi_data_out_r_39__N_2015[1] ;
    input resetn_c;
    input GND_net;
    input clk_enable_518;
    input n29080;
    input n26938;
    
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire [1:0]sync /* synthesis ASYNC_REG="TRUE" */ ;   // c:/s_links/sources/quad_decoder.v(106[30:34])
    wire [1:0]AB /* synthesis ASYNC_REG="TRUE" */ ;   // c:/s_links/sources/quad_decoder.v(106[36:38])
    wire \pin_intrpt[14]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[14] */ ;   // c:/s_links/sources/mcm_top.v(102[46:56])
    
    wire clk_1MHz_enable_213, n26211;
    wire [3:0]n2091;
    
    wire n28623;
    wire [31:0]quad_set;   // c:/s_links/sources/quad_decoder.v(40[31:39])
    
    wire n27, n19, n28942, n28941, n28935, n9746, n26747, quad_set_valid, 
        n9750, n29327, n29328, n11467;
    wire [31:0]n6106;
    
    wire n26955, n27094, n25843, n25845, n25863, n25865, n25883, 
        n25885, n25903, n25905, n25923, n25925, n25943, n25945, 
        n25963, n25965, n25983, n25985, n26003, n26005, n26023, 
        n26025, n26051, n26053, n26077, n26079, n26097, n26099, 
        n26125, n26127, n26157, n26159, n26205, n25170, n25169, 
        n25168, n25167, n25166, n25165, n25164, n25163, n25162, 
        n25161, n25160, n25159, n25158, n25157, n25156, n25155;
    
    FD1P3AX quad_count_i0_i0 (.D(n26211), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_2015[0] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX sync_i0 (.D(\quad_b[4] ), .CK(clk_1MHz), .Q(sync[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam sync_i0.GSR = "DISABLED";
    FD1S3AX AB_i0 (.D(sync[0]), .CK(clk_1MHz), .Q(AB[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam AB_i0.GSR = "DISABLED";
    FD1S3AX quad_buffer_i0 (.D(quad_count[0]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i0.GSR = "DISABLED";
    FD1S3JX state_FSM_i0 (.D(n28623), .CK(clk_1MHz), .PD(n29239), .Q(n2091[0]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i0.GSR = "DISABLED";
    FD1P3IX quad_set__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i0.GSR = "DISABLED";
    FD1P3IX quad_homing__i0 (.D(n29762), .SP(clk_enable_77), .CD(n29239), 
            .CK(clk), .Q(quad_homing[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam quad_homing__i0.GSR = "DISABLED";
    FD1P3IX quad_homing__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_77), .CD(n29239), 
            .CK(clk), .Q(quad_homing[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam quad_homing__i1.GSR = "DISABLED";
    FD1P3IX quad_set__i31 (.D(\spi_data_r[31] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i31.GSR = "DISABLED";
    FD1P3IX quad_set__i30 (.D(\spi_data_r[30] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i30.GSR = "DISABLED";
    FD1P3IX quad_set__i29 (.D(\spi_data_r[29] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i29.GSR = "DISABLED";
    FD1P3IX quad_set__i28 (.D(\spi_data_r[28] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i28.GSR = "DISABLED";
    FD1P3IX quad_set__i27 (.D(\spi_data_r[27] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i27.GSR = "DISABLED";
    FD1P3IX quad_set__i26 (.D(\spi_data_r[26] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i26.GSR = "DISABLED";
    FD1P3IX quad_set__i25 (.D(\spi_data_r[25] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i25.GSR = "DISABLED";
    FD1P3IX quad_set__i24 (.D(\spi_data_r[24] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i24.GSR = "DISABLED";
    FD1P3IX quad_set__i23 (.D(\spi_data_r[23] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i23.GSR = "DISABLED";
    FD1P3IX quad_set__i22 (.D(\spi_data_r[22] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i22.GSR = "DISABLED";
    FD1P3IX quad_set__i21 (.D(\spi_data_r[21] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i21.GSR = "DISABLED";
    FD1P3IX quad_set__i20 (.D(\spi_data_r[20] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i20.GSR = "DISABLED";
    FD1P3IX quad_set__i19 (.D(\spi_data_r[19] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i19.GSR = "DISABLED";
    FD1P3IX quad_set__i18 (.D(\spi_data_r[18] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i18.GSR = "DISABLED";
    FD1P3IX quad_set__i17 (.D(\spi_data_r[17] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i17.GSR = "DISABLED";
    FD1P3IX quad_set__i16 (.D(\spi_data_r[16] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i16.GSR = "DISABLED";
    FD1P3IX quad_set__i15 (.D(\spi_data_r[15] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i15.GSR = "DISABLED";
    FD1P3IX quad_set__i14 (.D(\spi_data_r[14] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i14.GSR = "DISABLED";
    FD1P3IX quad_set__i13 (.D(\spi_data_r[13] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i13.GSR = "DISABLED";
    FD1P3IX quad_set__i12 (.D(\spi_data_r[12] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i12.GSR = "DISABLED";
    FD1P3IX quad_set__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i11.GSR = "DISABLED";
    FD1P3IX quad_set__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i10.GSR = "DISABLED";
    FD1P3IX quad_set__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i9.GSR = "DISABLED";
    FD1P3IX quad_set__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i8.GSR = "DISABLED";
    FD1P3IX quad_set__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i7.GSR = "DISABLED";
    FD1P3IX quad_set__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i6.GSR = "DISABLED";
    FD1P3IX quad_set__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i5.GSR = "DISABLED";
    FD1P3IX quad_set__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i4.GSR = "DISABLED";
    FD1P3IX quad_set__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i3.GSR = "DISABLED";
    FD1P3IX quad_set__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i2.GSR = "DISABLED";
    FD1P3IX quad_set__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_162), .CD(n29239), 
            .CK(clk), .Q(quad_set[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i1.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(n2091[2]), .B(n2091[1]), .C(n2091[3]), .D(n27), 
         .Z(n19)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i1_4_lut.init = 16'hf10e;
    LUT4 i24_2_lut (.A(AB[1]), .B(AB[0]), .Z(n27)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam i24_2_lut.init = 16'h6666;
    FD1S3IX state_FSM_i3 (.D(n28942), .CK(clk_1MHz), .CD(n29239), .Q(n2091[3]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i3.GSR = "DISABLED";
    FD1S3IX state_FSM_i2 (.D(n28941), .CK(clk_1MHz), .CD(n29239), .Q(n2091[2]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i2.GSR = "DISABLED";
    FD1S3IX state_FSM_i1 (.D(n28935), .CK(clk_1MHz), .CD(n29239), .Q(n2091[1]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i1.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut (.A(n2091[3]), .B(AB[1]), .C(AB[0]), .D(n9746), 
         .Z(n26747)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i1_4_lut_4_lut.init = 16'h96c3;
    FD1S3IX quad_set_complete_451 (.D(quad_set_valid), .CK(clk_1MHz), .CD(n29239), 
            .Q(quad_set_complete)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_set_complete_451.GSR = "DISABLED";
    LUT4 AB_1__bdd_4_lut_23118 (.A(AB[1]), .B(n2091[1]), .C(AB[0]), .D(n9750), 
         .Z(n28935)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B (C (D))))) */ ;
    defparam AB_1__bdd_4_lut_23118.init = 16'h5848;
    FD1S3IX i41_407 (.D(spi_data_out_r_39__N_2098), .CK(clk), .CD(n29239), 
            .Q(spi_data_out_r_39__N_1910)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam i41_407.GSR = "DISABLED";
    LUT4 AB_1__bdd_4_lut (.A(AB[1]), .B(n2091[3]), .C(AB[0]), .D(n9746), 
         .Z(n28942)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam AB_1__bdd_4_lut.init = 16'ha484;
    LUT4 AB_1__bdd_4_lut_23119 (.A(AB[1]), .B(n2091[2]), .C(n9750), .D(AB[0]), 
         .Z(n28941)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B (D)))) */ ;
    defparam AB_1__bdd_4_lut_23119.init = 16'h44a8;
    PFUMX i23160 (.BLUT(n29327), .ALUT(n29328), .C0(AB[0]), .Z(n11467));
    LUT4 i33_4_lut_else_4_lut (.A(n2091[2]), .B(n2091[3]), .C(AB[1]), 
         .Z(n29327)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C)))) */ ;
    defparam i33_4_lut_else_4_lut.init = 16'h3d3d;
    LUT4 reduce_or_553_i1_2_lut (.A(n2091[3]), .B(n2091[0]), .Z(n9750)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam reduce_or_553_i1_2_lut.init = 16'heeee;
    LUT4 i33_4_lut (.A(n6106[31]), .B(quad_set[31]), .C(n26955), .D(n27094), 
         .Z(n25843)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut.init = 16'hac0c;
    LUT4 i33_4_lut_adj_840 (.A(n6106[30]), .B(quad_set[30]), .C(n26955), 
         .D(n27094), .Z(n25845)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_840.init = 16'hac0c;
    LUT4 i33_4_lut_adj_841 (.A(n6106[29]), .B(quad_set[29]), .C(n26955), 
         .D(n27094), .Z(n25863)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_841.init = 16'hac0c;
    LUT4 i33_4_lut_adj_842 (.A(n6106[28]), .B(quad_set[28]), .C(n26955), 
         .D(n27094), .Z(n25865)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_842.init = 16'hac0c;
    LUT4 i33_4_lut_adj_843 (.A(n6106[27]), .B(quad_set[27]), .C(n26955), 
         .D(n27094), .Z(n25883)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_843.init = 16'hac0c;
    LUT4 i33_4_lut_adj_844 (.A(n6106[26]), .B(quad_set[26]), .C(n26955), 
         .D(n27094), .Z(n25885)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_844.init = 16'hac0c;
    LUT4 i33_4_lut_adj_845 (.A(n6106[25]), .B(quad_set[25]), .C(n26955), 
         .D(n27094), .Z(n25903)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_845.init = 16'hac0c;
    LUT4 i33_4_lut_adj_846 (.A(n6106[24]), .B(quad_set[24]), .C(n26955), 
         .D(n27094), .Z(n25905)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_846.init = 16'hac0c;
    LUT4 i33_4_lut_adj_847 (.A(n6106[23]), .B(quad_set[23]), .C(n26955), 
         .D(n27094), .Z(n25923)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_847.init = 16'hac0c;
    LUT4 i33_4_lut_adj_848 (.A(n6106[22]), .B(quad_set[22]), .C(n26955), 
         .D(n27094), .Z(n25925)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_848.init = 16'hac0c;
    LUT4 i33_4_lut_adj_849 (.A(n6106[21]), .B(quad_set[21]), .C(n26955), 
         .D(n27094), .Z(n25943)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_849.init = 16'hac0c;
    LUT4 i33_4_lut_adj_850 (.A(n6106[20]), .B(quad_set[20]), .C(n26955), 
         .D(n27094), .Z(n25945)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_850.init = 16'hac0c;
    LUT4 i33_4_lut_adj_851 (.A(n6106[19]), .B(quad_set[19]), .C(n26955), 
         .D(n27094), .Z(n25963)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_851.init = 16'hac0c;
    LUT4 i33_4_lut_adj_852 (.A(n6106[18]), .B(quad_set[18]), .C(n26955), 
         .D(n27094), .Z(n25965)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_852.init = 16'hac0c;
    LUT4 i33_4_lut_adj_853 (.A(n6106[17]), .B(quad_set[17]), .C(n26955), 
         .D(n27094), .Z(n25983)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_853.init = 16'hac0c;
    LUT4 i33_4_lut_adj_854 (.A(n6106[16]), .B(quad_set[16]), .C(n26955), 
         .D(n27094), .Z(n25985)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_854.init = 16'hac0c;
    LUT4 i33_4_lut_adj_855 (.A(n6106[15]), .B(quad_set[15]), .C(n26955), 
         .D(n27094), .Z(n26003)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_855.init = 16'hac0c;
    LUT4 i33_4_lut_adj_856 (.A(n6106[14]), .B(quad_set[14]), .C(n26955), 
         .D(n27094), .Z(n26005)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_856.init = 16'hac0c;
    LUT4 i33_4_lut_adj_857 (.A(n6106[13]), .B(quad_set[13]), .C(n26955), 
         .D(n27094), .Z(n26023)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_857.init = 16'hac0c;
    LUT4 i33_4_lut_adj_858 (.A(n6106[12]), .B(quad_set[12]), .C(n26955), 
         .D(n27094), .Z(n26025)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_858.init = 16'hac0c;
    LUT4 i33_4_lut_adj_859 (.A(n6106[11]), .B(quad_set[11]), .C(n26955), 
         .D(n27094), .Z(n26051)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_859.init = 16'hac0c;
    LUT4 i33_4_lut_adj_860 (.A(n6106[10]), .B(quad_set[10]), .C(n26955), 
         .D(n27094), .Z(n26053)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_860.init = 16'hac0c;
    LUT4 i33_4_lut_adj_861 (.A(n6106[9]), .B(quad_set[9]), .C(n26955), 
         .D(n27094), .Z(n26077)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_861.init = 16'hac0c;
    LUT4 i33_4_lut_adj_862 (.A(n6106[8]), .B(quad_set[8]), .C(n26955), 
         .D(n27094), .Z(n26079)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_862.init = 16'hac0c;
    LUT4 i33_4_lut_adj_863 (.A(n6106[7]), .B(quad_set[7]), .C(n26955), 
         .D(n27094), .Z(n26097)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_863.init = 16'hac0c;
    LUT4 i33_4_lut_adj_864 (.A(n6106[6]), .B(quad_set[6]), .C(n26955), 
         .D(n27094), .Z(n26099)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_864.init = 16'hac0c;
    LUT4 i33_4_lut_adj_865 (.A(n6106[5]), .B(quad_set[5]), .C(n26955), 
         .D(n27094), .Z(n26125)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_865.init = 16'hac0c;
    LUT4 i33_4_lut_adj_866 (.A(n6106[4]), .B(quad_set[4]), .C(n26955), 
         .D(n27094), .Z(n26127)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_866.init = 16'hac0c;
    LUT4 i33_4_lut_adj_867 (.A(n6106[3]), .B(quad_set[3]), .C(n26955), 
         .D(n27094), .Z(n26157)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_867.init = 16'hac0c;
    FD1S3AX quad_buffer_i31 (.D(quad_count[31]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i31.GSR = "DISABLED";
    FD1S3AX quad_buffer_i30 (.D(quad_count[30]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i30.GSR = "DISABLED";
    FD1S3AX quad_buffer_i29 (.D(quad_count[29]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i29.GSR = "DISABLED";
    FD1S3AX quad_buffer_i28 (.D(quad_count[28]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i28.GSR = "DISABLED";
    FD1S3AX quad_buffer_i27 (.D(quad_count[27]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i27.GSR = "DISABLED";
    FD1S3AX quad_buffer_i26 (.D(quad_count[26]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i26.GSR = "DISABLED";
    FD1S3AX quad_buffer_i25 (.D(quad_count[25]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i25.GSR = "DISABLED";
    FD1S3AX quad_buffer_i24 (.D(quad_count[24]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i24.GSR = "DISABLED";
    FD1S3AX quad_buffer_i23 (.D(quad_count[23]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i23.GSR = "DISABLED";
    FD1S3AX quad_buffer_i22 (.D(quad_count[22]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i22.GSR = "DISABLED";
    FD1S3AX quad_buffer_i21 (.D(quad_count[21]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i21.GSR = "DISABLED";
    FD1S3AX quad_buffer_i20 (.D(quad_count[20]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i20.GSR = "DISABLED";
    FD1S3AX quad_buffer_i19 (.D(quad_count[19]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i19.GSR = "DISABLED";
    FD1S3AX quad_buffer_i18 (.D(quad_count[18]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i18.GSR = "DISABLED";
    FD1S3AX quad_buffer_i17 (.D(quad_count[17]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i17.GSR = "DISABLED";
    LUT4 i33_4_lut_adj_868 (.A(n6106[2]), .B(quad_set[2]), .C(n26955), 
         .D(n27094), .Z(n26159)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_868.init = 16'hac0c;
    LUT4 i33_4_lut_adj_869 (.A(n6106[1]), .B(quad_set[1]), .C(n26955), 
         .D(n27094), .Z(n26205)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_869.init = 16'hac0c;
    FD1S3AX quad_buffer_i16 (.D(quad_count[16]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i16.GSR = "DISABLED";
    FD1S3AX quad_buffer_i15 (.D(quad_count[15]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i15.GSR = "DISABLED";
    FD1S3AX quad_buffer_i14 (.D(quad_count[14]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i14.GSR = "DISABLED";
    FD1S3AX quad_buffer_i13 (.D(quad_count[13]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i13.GSR = "DISABLED";
    FD1S3AX quad_buffer_i12 (.D(quad_count[12]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i12.GSR = "DISABLED";
    FD1S3AX quad_buffer_i11 (.D(quad_count[11]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i11.GSR = "DISABLED";
    FD1S3AX quad_buffer_i10 (.D(quad_count[10]), .CK(\pin_intrpt[14] ), 
            .Q(quad_buffer[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i10.GSR = "DISABLED";
    FD1S3AX quad_buffer_i9 (.D(quad_count[9]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i9.GSR = "DISABLED";
    FD1S3AX quad_buffer_i8 (.D(quad_count[8]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i8.GSR = "DISABLED";
    FD1S3AX quad_buffer_i7 (.D(quad_count[7]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i7.GSR = "DISABLED";
    FD1S3AX quad_buffer_i6 (.D(quad_count[6]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i6.GSR = "DISABLED";
    FD1S3AX quad_buffer_i5 (.D(quad_count[5]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i5.GSR = "DISABLED";
    FD1S3AX quad_buffer_i4 (.D(quad_count[4]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i4.GSR = "DISABLED";
    FD1S3AX quad_buffer_i3 (.D(quad_count[3]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i3.GSR = "DISABLED";
    FD1S3AX quad_buffer_i2 (.D(quad_count[2]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i2.GSR = "DISABLED";
    FD1S3AX quad_buffer_i1 (.D(quad_count[1]), .CK(\pin_intrpt[14] ), .Q(quad_buffer[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i1.GSR = "DISABLED";
    FD1S3AX AB_i1 (.D(sync[1]), .CK(clk_1MHz), .Q(AB[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam AB_i1.GSR = "DISABLED";
    FD1S3AX sync_i1 (.D(\quad_a[4] ), .CK(clk_1MHz), .Q(sync[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam sync_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_2015[31] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i31 (.D(\spi_data_out_r_39__N_2015[30] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i30 (.D(\spi_data_out_r_39__N_2015[29] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i29 (.D(\spi_data_out_r_39__N_2015[28] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i28 (.D(\spi_data_out_r_39__N_2015[27] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i27 (.D(\spi_data_out_r_39__N_2015[26] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i26 (.D(\spi_data_out_r_39__N_2015[25] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i25 (.D(\spi_data_out_r_39__N_2015[24] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i24 (.D(\spi_data_out_r_39__N_2015[23] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i23 (.D(\spi_data_out_r_39__N_2015[22] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i22 (.D(\spi_data_out_r_39__N_2015[21] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i21 (.D(\spi_data_out_r_39__N_2015[20] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i20 (.D(\spi_data_out_r_39__N_2015[19] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i19 (.D(\spi_data_out_r_39__N_2015[18] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i18 (.D(\spi_data_out_r_39__N_2015[17] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i17 (.D(\spi_data_out_r_39__N_2015[16] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i16 (.D(\spi_data_out_r_39__N_2015[15] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_2015[14] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_2015[13] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_2015[12] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_2015[11] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_2015[10] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_2015[9] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_2015[8] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_2015[7] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_2015[6] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_2015[5] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_2015[4] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_2015[3] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_2015[2] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_2015[1] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1870[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    LUT4 i33_4_lut_then_4_lut (.A(n2091[2]), .B(n2091[3]), .C(AB[1]), 
         .D(n2091[1]), .Z(n29328)) /* synthesis lut_function=(A+(B+!(C (D)+!C !(D)))) */ ;
    defparam i33_4_lut_then_4_lut.init = 16'heffe;
    LUT4 reduce_or_558_i1_2_lut (.A(n2091[2]), .B(n2091[1]), .Z(n9746)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam reduce_or_558_i1_2_lut.init = 16'heeee;
    FD1P3AX quad_count_i0_i31 (.D(n25843), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i31.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i30 (.D(n25845), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i30.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i29 (.D(n25863), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i29.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i28 (.D(n25865), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i28.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i27 (.D(n25883), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i27.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i26 (.D(n25885), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i26.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i25 (.D(n25903), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i25.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i24 (.D(n25905), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i24.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i23 (.D(n25923), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i23.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i22 (.D(n25925), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i22.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i21 (.D(n25943), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i21.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i20 (.D(n25945), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i20.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i19 (.D(n25963), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i19.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i18 (.D(n25965), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i18.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i17 (.D(n25983), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i17.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i16 (.D(n25985), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i16.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i15 (.D(n26003), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i15.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i14 (.D(n26005), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i14.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i13 (.D(n26023), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i13.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i12 (.D(n26025), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i12.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i11 (.D(n26051), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i11.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i10 (.D(n26053), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i10.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i9 (.D(n26077), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i9.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i8 (.D(n26079), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i8.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i7 (.D(n26097), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i7.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i6 (.D(n26099), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i6.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i5 (.D(n26125), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i5.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i4 (.D(n26127), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i4.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i3 (.D(n26157), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i3.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i2 (.D(n26159), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i1 (.D(n26205), .SP(clk_1MHz_enable_213), .CK(clk_1MHz), 
            .Q(quad_count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i1.GSR = "DISABLED";
    CCU2D add_1947_33 (.A0(resetn_c), .B0(n11467), .C0(quad_count[30]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[31]), 
          .D1(GND_net), .CIN(n25170), .S0(n6106[30]), .S1(n6106[31]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_33.INIT0 = 16'hd2d2;
    defparam add_1947_33.INIT1 = 16'hd2d2;
    defparam add_1947_33.INJECT1_0 = "NO";
    defparam add_1947_33.INJECT1_1 = "NO";
    CCU2D add_1947_31 (.A0(resetn_c), .B0(n11467), .C0(quad_count[28]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[29]), 
          .D1(GND_net), .CIN(n25169), .COUT(n25170), .S0(n6106[28]), 
          .S1(n6106[29]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_31.INIT0 = 16'hd2d2;
    defparam add_1947_31.INIT1 = 16'hd2d2;
    defparam add_1947_31.INJECT1_0 = "NO";
    defparam add_1947_31.INJECT1_1 = "NO";
    CCU2D add_1947_29 (.A0(resetn_c), .B0(n11467), .C0(quad_count[26]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[27]), 
          .D1(GND_net), .CIN(n25168), .COUT(n25169), .S0(n6106[26]), 
          .S1(n6106[27]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_29.INIT0 = 16'hd2d2;
    defparam add_1947_29.INIT1 = 16'hd2d2;
    defparam add_1947_29.INJECT1_0 = "NO";
    defparam add_1947_29.INJECT1_1 = "NO";
    CCU2D add_1947_27 (.A0(resetn_c), .B0(n11467), .C0(quad_count[24]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[25]), 
          .D1(GND_net), .CIN(n25167), .COUT(n25168), .S0(n6106[24]), 
          .S1(n6106[25]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_27.INIT0 = 16'hd2d2;
    defparam add_1947_27.INIT1 = 16'hd2d2;
    defparam add_1947_27.INJECT1_0 = "NO";
    defparam add_1947_27.INJECT1_1 = "NO";
    CCU2D add_1947_25 (.A0(resetn_c), .B0(n11467), .C0(quad_count[22]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[23]), 
          .D1(GND_net), .CIN(n25166), .COUT(n25167), .S0(n6106[22]), 
          .S1(n6106[23]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_25.INIT0 = 16'hd2d2;
    defparam add_1947_25.INIT1 = 16'hd2d2;
    defparam add_1947_25.INJECT1_0 = "NO";
    defparam add_1947_25.INJECT1_1 = "NO";
    CCU2D add_1947_23 (.A0(resetn_c), .B0(n11467), .C0(quad_count[20]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[21]), 
          .D1(GND_net), .CIN(n25165), .COUT(n25166), .S0(n6106[20]), 
          .S1(n6106[21]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_23.INIT0 = 16'hd2d2;
    defparam add_1947_23.INIT1 = 16'hd2d2;
    defparam add_1947_23.INJECT1_0 = "NO";
    defparam add_1947_23.INJECT1_1 = "NO";
    LUT4 AB_1__bdd_4_lut_23114 (.A(AB[1]), .B(n2091[0]), .C(AB[0]), .D(n9746), 
         .Z(n28623)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B (C+!(D)))) */ ;
    defparam AB_1__bdd_4_lut_23114.init = 16'h8584;
    CCU2D add_1947_21 (.A0(resetn_c), .B0(n11467), .C0(quad_count[18]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[19]), 
          .D1(GND_net), .CIN(n25164), .COUT(n25165), .S0(n6106[18]), 
          .S1(n6106[19]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_21.INIT0 = 16'hd2d2;
    defparam add_1947_21.INIT1 = 16'hd2d2;
    defparam add_1947_21.INJECT1_0 = "NO";
    defparam add_1947_21.INJECT1_1 = "NO";
    CCU2D add_1947_19 (.A0(resetn_c), .B0(n11467), .C0(quad_count[16]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[17]), 
          .D1(GND_net), .CIN(n25163), .COUT(n25164), .S0(n6106[16]), 
          .S1(n6106[17]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_19.INIT0 = 16'hd2d2;
    defparam add_1947_19.INIT1 = 16'hd2d2;
    defparam add_1947_19.INJECT1_0 = "NO";
    defparam add_1947_19.INJECT1_1 = "NO";
    CCU2D add_1947_17 (.A0(resetn_c), .B0(n11467), .C0(quad_count[14]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[15]), 
          .D1(GND_net), .CIN(n25162), .COUT(n25163), .S0(n6106[14]), 
          .S1(n6106[15]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_17.INIT0 = 16'hd2d2;
    defparam add_1947_17.INIT1 = 16'hd2d2;
    defparam add_1947_17.INJECT1_0 = "NO";
    defparam add_1947_17.INJECT1_1 = "NO";
    CCU2D add_1947_15 (.A0(resetn_c), .B0(n11467), .C0(quad_count[12]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[13]), 
          .D1(GND_net), .CIN(n25161), .COUT(n25162), .S0(n6106[12]), 
          .S1(n6106[13]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_15.INIT0 = 16'hd2d2;
    defparam add_1947_15.INIT1 = 16'hd2d2;
    defparam add_1947_15.INJECT1_0 = "NO";
    defparam add_1947_15.INJECT1_1 = "NO";
    CCU2D add_1947_13 (.A0(resetn_c), .B0(n11467), .C0(quad_count[10]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[11]), 
          .D1(GND_net), .CIN(n25160), .COUT(n25161), .S0(n6106[10]), 
          .S1(n6106[11]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_13.INIT0 = 16'hd2d2;
    defparam add_1947_13.INIT1 = 16'hd2d2;
    defparam add_1947_13.INJECT1_0 = "NO";
    defparam add_1947_13.INJECT1_1 = "NO";
    CCU2D add_1947_11 (.A0(resetn_c), .B0(n11467), .C0(quad_count[8]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[9]), 
          .D1(GND_net), .CIN(n25159), .COUT(n25160), .S0(n6106[8]), 
          .S1(n6106[9]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_11.INIT0 = 16'hd2d2;
    defparam add_1947_11.INIT1 = 16'hd2d2;
    defparam add_1947_11.INJECT1_0 = "NO";
    defparam add_1947_11.INJECT1_1 = "NO";
    CCU2D add_1947_9 (.A0(resetn_c), .B0(n11467), .C0(quad_count[6]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[7]), 
          .D1(GND_net), .CIN(n25158), .COUT(n25159), .S0(n6106[6]), 
          .S1(n6106[7]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_9.INIT0 = 16'hd2d2;
    defparam add_1947_9.INIT1 = 16'hd2d2;
    defparam add_1947_9.INJECT1_0 = "NO";
    defparam add_1947_9.INJECT1_1 = "NO";
    CCU2D add_1947_7 (.A0(resetn_c), .B0(n11467), .C0(quad_count[4]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[5]), 
          .D1(GND_net), .CIN(n25157), .COUT(n25158), .S0(n6106[4]), 
          .S1(n6106[5]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_7.INIT0 = 16'hd2d2;
    defparam add_1947_7.INIT1 = 16'hd2d2;
    defparam add_1947_7.INJECT1_0 = "NO";
    defparam add_1947_7.INJECT1_1 = "NO";
    CCU2D add_1947_5 (.A0(resetn_c), .B0(n11467), .C0(quad_count[2]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[3]), 
          .D1(GND_net), .CIN(n25156), .COUT(n25157), .S0(n6106[2]), 
          .S1(n6106[3]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_5.INIT0 = 16'hd2d2;
    defparam add_1947_5.INIT1 = 16'hd2d2;
    defparam add_1947_5.INJECT1_0 = "NO";
    defparam add_1947_5.INJECT1_1 = "NO";
    CCU2D add_1947_3 (.A0(resetn_c), .B0(n11467), .C0(quad_count[0]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11467), .C1(quad_count[1]), 
          .D1(GND_net), .CIN(n25155), .COUT(n25156), .S0(n6106[0]), 
          .S1(n6106[1]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_3.INIT0 = 16'h2d2d;
    defparam add_1947_3.INIT1 = 16'hd2d2;
    defparam add_1947_3.INJECT1_0 = "NO";
    defparam add_1947_3.INJECT1_1 = "NO";
    CCU2D add_1947_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(resetn_c), .B1(n11467), .C1(GND_net), .D1(GND_net), .COUT(n25155));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1947_1.INIT0 = 16'hF000;
    defparam add_1947_1.INIT1 = 16'hdddd;
    defparam add_1947_1.INJECT1_0 = "NO";
    defparam add_1947_1.INJECT1_1 = "NO";
    FD1P3IX quad_set_valid_404 (.D(n29080), .SP(clk_enable_518), .CD(n29239), 
            .CK(clk), .Q(quad_set_valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set_valid_404.GSR = "DISABLED";
    LUT4 i22885_4_lut (.A(resetn_c), .B(quad_set_valid), .C(n26747), .D(n26938), 
         .Z(clk_1MHz_enable_213)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i22885_4_lut.init = 16'hffdf;
    LUT4 i33_4_lut_adj_870 (.A(n6106[0]), .B(quad_set[0]), .C(n26955), 
         .D(n27094), .Z(n26211)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i33_4_lut_adj_870.init = 16'hac0c;
    LUT4 i2_4_lut (.A(n26938), .B(resetn_c), .C(n19), .D(quad_set_valid), 
         .Z(n26955)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;
    defparam i2_4_lut.init = 16'hfbff;
    LUT4 i1_3_lut (.A(resetn_c), .B(n26938), .C(n19), .Z(n27094)) /* synthesis lut_function=(A ((C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i1_3_lut.init = 16'ha2a2;
    
endmodule
//
// Verilog Description of module \quad_decoder(DEV_ID=1) 
//

module \quad_decoder(DEV_ID=1)  (clk, clk_enable_286, n29239, n29762, 
            quad_count, clk_1MHz, \spi_data_out_r_39__N_1168[0] , \spi_data_out_r_39__N_1313[0] , 
            \quad_b[1] , quad_buffer, \pin_intrpt[5] , clk_enable_467, 
            \spi_data_r[0] , quad_set_complete, spi_data_out_r_39__N_1208, 
            spi_data_out_r_39__N_1396, resetn_c, GND_net, \quad_a[1] , 
            \spi_data_out_r_39__N_1168[31] , \spi_data_out_r_39__N_1313[31] , 
            \spi_data_out_r_39__N_1168[30] , \spi_data_out_r_39__N_1313[30] , 
            \spi_data_out_r_39__N_1168[29] , \spi_data_out_r_39__N_1313[29] , 
            \spi_data_out_r_39__N_1168[28] , \spi_data_out_r_39__N_1313[28] , 
            \spi_data_out_r_39__N_1168[27] , \spi_data_out_r_39__N_1313[27] , 
            \spi_data_out_r_39__N_1168[26] , \spi_data_out_r_39__N_1313[26] , 
            \spi_data_out_r_39__N_1168[25] , \spi_data_out_r_39__N_1313[25] , 
            \spi_data_out_r_39__N_1168[24] , \spi_data_out_r_39__N_1313[24] , 
            \spi_data_out_r_39__N_1168[23] , \spi_data_out_r_39__N_1313[23] , 
            \spi_data_out_r_39__N_1168[22] , \spi_data_out_r_39__N_1313[22] , 
            \spi_data_out_r_39__N_1168[21] , \spi_data_out_r_39__N_1313[21] , 
            \spi_data_out_r_39__N_1168[20] , \spi_data_out_r_39__N_1313[20] , 
            \spi_data_out_r_39__N_1168[19] , \spi_data_out_r_39__N_1313[19] , 
            \spi_data_out_r_39__N_1168[18] , \spi_data_out_r_39__N_1313[18] , 
            \spi_data_out_r_39__N_1168[17] , \spi_data_out_r_39__N_1313[17] , 
            \spi_data_out_r_39__N_1168[16] , \spi_data_out_r_39__N_1313[16] , 
            \spi_data_out_r_39__N_1168[15] , \spi_data_out_r_39__N_1313[15] , 
            \spi_data_out_r_39__N_1168[14] , \spi_data_out_r_39__N_1313[14] , 
            \spi_data_out_r_39__N_1168[13] , \spi_data_out_r_39__N_1313[13] , 
            \spi_data_out_r_39__N_1168[12] , \spi_data_out_r_39__N_1313[12] , 
            \spi_data_out_r_39__N_1168[11] , \spi_data_out_r_39__N_1313[11] , 
            \spi_data_out_r_39__N_1168[10] , \spi_data_out_r_39__N_1313[10] , 
            \spi_data_out_r_39__N_1168[9] , \spi_data_out_r_39__N_1313[9] , 
            \spi_data_out_r_39__N_1168[8] , \spi_data_out_r_39__N_1313[8] , 
            \spi_data_out_r_39__N_1168[7] , \spi_data_out_r_39__N_1313[7] , 
            \spi_data_out_r_39__N_1168[6] , \spi_data_out_r_39__N_1313[6] , 
            \spi_data_out_r_39__N_1168[5] , \spi_data_out_r_39__N_1313[5] , 
            \spi_data_out_r_39__N_1168[4] , \spi_data_out_r_39__N_1313[4] , 
            \spi_data_out_r_39__N_1168[3] , \spi_data_out_r_39__N_1313[3] , 
            \spi_data_out_r_39__N_1168[2] , \spi_data_out_r_39__N_1313[2] , 
            \spi_data_out_r_39__N_1168[1] , \spi_data_out_r_39__N_1313[1] , 
            \quad_homing[1] , \spi_data_r[1] , \spi_data_r[2] , \spi_data_r[3] , 
            \spi_data_r[4] , \spi_data_r[5] , \spi_data_r[6] , \spi_data_r[7] , 
            \spi_data_r[8] , \spi_data_r[9] , \spi_data_r[10] , \spi_data_r[11] , 
            \spi_data_r[12] , \spi_data_r[13] , \spi_data_r[14] , \spi_data_r[15] , 
            \spi_data_r[16] , \spi_data_r[17] , \spi_data_r[18] , \spi_data_r[19] , 
            \spi_data_r[20] , \spi_data_r[21] , \spi_data_r[22] , \spi_data_r[23] , 
            \spi_data_r[24] , \spi_data_r[25] , \spi_data_r[26] , \spi_data_r[27] , 
            \spi_data_r[28] , \spi_data_r[29] , \spi_data_r[30] , \spi_data_r[31] , 
            clk_enable_502, n29084, n12716, n26963, pin_io_out_14, 
            n27636) /* synthesis syn_module_defined=1 */ ;
    input clk;
    input clk_enable_286;
    input n29239;
    input n29762;
    output [31:0]quad_count;
    input clk_1MHz;
    output \spi_data_out_r_39__N_1168[0] ;
    input \spi_data_out_r_39__N_1313[0] ;
    input \quad_b[1] ;
    output [31:0]quad_buffer;
    input \pin_intrpt[5] ;
    input clk_enable_467;
    input \spi_data_r[0] ;
    output quad_set_complete;
    output spi_data_out_r_39__N_1208;
    input spi_data_out_r_39__N_1396;
    input resetn_c;
    input GND_net;
    input \quad_a[1] ;
    output \spi_data_out_r_39__N_1168[31] ;
    input \spi_data_out_r_39__N_1313[31] ;
    output \spi_data_out_r_39__N_1168[30] ;
    input \spi_data_out_r_39__N_1313[30] ;
    output \spi_data_out_r_39__N_1168[29] ;
    input \spi_data_out_r_39__N_1313[29] ;
    output \spi_data_out_r_39__N_1168[28] ;
    input \spi_data_out_r_39__N_1313[28] ;
    output \spi_data_out_r_39__N_1168[27] ;
    input \spi_data_out_r_39__N_1313[27] ;
    output \spi_data_out_r_39__N_1168[26] ;
    input \spi_data_out_r_39__N_1313[26] ;
    output \spi_data_out_r_39__N_1168[25] ;
    input \spi_data_out_r_39__N_1313[25] ;
    output \spi_data_out_r_39__N_1168[24] ;
    input \spi_data_out_r_39__N_1313[24] ;
    output \spi_data_out_r_39__N_1168[23] ;
    input \spi_data_out_r_39__N_1313[23] ;
    output \spi_data_out_r_39__N_1168[22] ;
    input \spi_data_out_r_39__N_1313[22] ;
    output \spi_data_out_r_39__N_1168[21] ;
    input \spi_data_out_r_39__N_1313[21] ;
    output \spi_data_out_r_39__N_1168[20] ;
    input \spi_data_out_r_39__N_1313[20] ;
    output \spi_data_out_r_39__N_1168[19] ;
    input \spi_data_out_r_39__N_1313[19] ;
    output \spi_data_out_r_39__N_1168[18] ;
    input \spi_data_out_r_39__N_1313[18] ;
    output \spi_data_out_r_39__N_1168[17] ;
    input \spi_data_out_r_39__N_1313[17] ;
    output \spi_data_out_r_39__N_1168[16] ;
    input \spi_data_out_r_39__N_1313[16] ;
    output \spi_data_out_r_39__N_1168[15] ;
    input \spi_data_out_r_39__N_1313[15] ;
    output \spi_data_out_r_39__N_1168[14] ;
    input \spi_data_out_r_39__N_1313[14] ;
    output \spi_data_out_r_39__N_1168[13] ;
    input \spi_data_out_r_39__N_1313[13] ;
    output \spi_data_out_r_39__N_1168[12] ;
    input \spi_data_out_r_39__N_1313[12] ;
    output \spi_data_out_r_39__N_1168[11] ;
    input \spi_data_out_r_39__N_1313[11] ;
    output \spi_data_out_r_39__N_1168[10] ;
    input \spi_data_out_r_39__N_1313[10] ;
    output \spi_data_out_r_39__N_1168[9] ;
    input \spi_data_out_r_39__N_1313[9] ;
    output \spi_data_out_r_39__N_1168[8] ;
    input \spi_data_out_r_39__N_1313[8] ;
    output \spi_data_out_r_39__N_1168[7] ;
    input \spi_data_out_r_39__N_1313[7] ;
    output \spi_data_out_r_39__N_1168[6] ;
    input \spi_data_out_r_39__N_1313[6] ;
    output \spi_data_out_r_39__N_1168[5] ;
    input \spi_data_out_r_39__N_1313[5] ;
    output \spi_data_out_r_39__N_1168[4] ;
    input \spi_data_out_r_39__N_1313[4] ;
    output \spi_data_out_r_39__N_1168[3] ;
    input \spi_data_out_r_39__N_1313[3] ;
    output \spi_data_out_r_39__N_1168[2] ;
    input \spi_data_out_r_39__N_1313[2] ;
    output \spi_data_out_r_39__N_1168[1] ;
    input \spi_data_out_r_39__N_1313[1] ;
    output \quad_homing[1] ;
    input \spi_data_r[1] ;
    input \spi_data_r[2] ;
    input \spi_data_r[3] ;
    input \spi_data_r[4] ;
    input \spi_data_r[5] ;
    input \spi_data_r[6] ;
    input \spi_data_r[7] ;
    input \spi_data_r[8] ;
    input \spi_data_r[9] ;
    input \spi_data_r[10] ;
    input \spi_data_r[11] ;
    input \spi_data_r[12] ;
    input \spi_data_r[13] ;
    input \spi_data_r[14] ;
    input \spi_data_r[15] ;
    input \spi_data_r[16] ;
    input \spi_data_r[17] ;
    input \spi_data_r[18] ;
    input \spi_data_r[19] ;
    input \spi_data_r[20] ;
    input \spi_data_r[21] ;
    input \spi_data_r[22] ;
    input \spi_data_r[23] ;
    input \spi_data_r[24] ;
    input \spi_data_r[25] ;
    input \spi_data_r[26] ;
    input \spi_data_r[27] ;
    input \spi_data_r[28] ;
    input \spi_data_r[29] ;
    input \spi_data_r[30] ;
    input \spi_data_r[31] ;
    input clk_enable_502;
    input n29084;
    input n12716;
    input n26963;
    input pin_io_out_14;
    output n27636;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire [1:0]sync /* synthesis ASYNC_REG="TRUE" */ ;   // c:/s_links/sources/quad_decoder.v(106[30:34])
    wire [1:0]AB /* synthesis ASYNC_REG="TRUE" */ ;   // c:/s_links/sources/quad_decoder.v(106[36:38])
    wire \pin_intrpt[5]  /* synthesis is_clock=1, SET_AS_NETWORK=pin_intrpt[5] */ ;   // c:/s_links/sources/mcm_top.v(102[46:56])
    wire [1:0]quad_homing;   // c:/s_links/sources/quad_decoder.v(41[19:30])
    
    wire clk_1MHz_enable_309, n26141;
    wire [3:0]n1521;
    
    wire n11361, n11558, n28864;
    wire [31:0]quad_set;   // c:/s_links/sources/quad_decoder.v(40[31:39])
    
    wire n6, n9488, n8, n26753, n28609, quad_set_valid, n28608, 
        n25090;
    wire [31:0]n6366;
    
    wire n25089, n25088, n25087, n25086, n25085, n25084, n25083, 
        n25082, n25081, n25080, n25079, n25078, n25077, n25076, 
        n25075, n25837, n25835, n25857, n25855, n25877, n25875, 
        n25897, n25895, n25917, n25915, n25937, n25935, n25957, 
        n25955, n25977, n25975, n25997, n25995, n26017, n26015, 
        n26037, n26035, n26065, n26063, n26091, n26089, n26111, 
        n26109, n26139, n26137, n26167, n3, n27061, n4, n12;
    
    FD1P3IX quad_homing__i0 (.D(n29762), .SP(clk_enable_286), .CD(n29239), 
            .CK(clk), .Q(quad_homing[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam quad_homing__i0.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i0 (.D(n26141), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_1313[0] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX sync_i0 (.D(\quad_b[1] ), .CK(clk_1MHz), .Q(sync[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam sync_i0.GSR = "DISABLED";
    FD1S3AX AB_i0 (.D(sync[0]), .CK(clk_1MHz), .Q(AB[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam AB_i0.GSR = "DISABLED";
    FD1S3AX quad_buffer_i0 (.D(quad_count[0]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i0.GSR = "DISABLED";
    LUT4 i5154_3_lut_4_lut (.A(AB[0]), .B(AB[1]), .C(n1521[3]), .D(n11361), 
         .Z(n11558)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // c:/s_links/sources/quad_decoder.v(162[19:30])
    defparam i5154_3_lut_4_lut.init = 16'hbfb0;
    FD1S3JX state_FSM_i0 (.D(n28864), .CK(clk_1MHz), .PD(n29239), .Q(n1521[0]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i0.GSR = "DISABLED";
    FD1P3IX quad_set__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i0.GSR = "DISABLED";
    LUT4 i4712_4_lut_4_lut (.A(n1521[2]), .B(AB[0]), .C(AB[1]), .D(n6), 
         .Z(n9488)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C (D))))) */ ;   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam i4712_4_lut_4_lut.init = 16'h3828;
    LUT4 i1_4_lut_4_lut (.A(n1521[3]), .B(AB[0]), .C(AB[1]), .D(n8), 
         .Z(n26753)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i1_4_lut_4_lut.init = 16'h96c3;
    LUT4 n8_bdd_4_lut_23098 (.A(n8), .B(n1521[3]), .C(AB[1]), .D(AB[0]), 
         .Z(n28609)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C (D)))+!A (B (C (D)+!C !(D)))) */ ;
    defparam n8_bdd_4_lut_23098.init = 16'he00c;
    LUT4 i5153_4_lut (.A(AB[0]), .B(AB[1]), .C(n1521[2]), .D(n1521[1]), 
         .Z(n11361)) /* synthesis lut_function=(A (B (C+!(D))+!B (C+(D)))+!A (B+!(C))) */ ;
    defparam i5153_4_lut.init = 16'he7ed;
    FD1S3IX quad_set_complete_451 (.D(quad_set_valid), .CK(clk_1MHz), .CD(n29239), 
            .Q(quad_set_complete)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_set_complete_451.GSR = "DISABLED";
    FD1S3IX i41_407 (.D(spi_data_out_r_39__N_1396), .CK(clk), .CD(n29239), 
            .Q(spi_data_out_r_39__N_1208)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam i41_407.GSR = "DISABLED";
    LUT4 n6_bdd_4_lut (.A(n6), .B(n1521[1]), .C(AB[0]), .D(AB[1]), .Z(n28608)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C (D)+!C !(D))+!B))) */ ;
    defparam n6_bdd_4_lut.init = 16'h0ce0;
    FD1S3IX state_FSM_i3 (.D(n28609), .CK(clk_1MHz), .CD(n29239), .Q(n1521[3]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i3.GSR = "DISABLED";
    FD1S3IX state_FSM_i2 (.D(n9488), .CK(clk_1MHz), .CD(n29239), .Q(n1521[2]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i2.GSR = "DISABLED";
    FD1S3IX state_FSM_i1 (.D(n28608), .CK(clk_1MHz), .CD(n29239), .Q(n1521[1]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i1.GSR = "DISABLED";
    CCU2D add_2079_33 (.A0(resetn_c), .B0(n11558), .C0(quad_count[30]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[31]), 
          .D1(GND_net), .CIN(n25090), .S0(n6366[30]), .S1(n6366[31]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_33.INIT0 = 16'hd2d2;
    defparam add_2079_33.INIT1 = 16'hd2d2;
    defparam add_2079_33.INJECT1_0 = "NO";
    defparam add_2079_33.INJECT1_1 = "NO";
    CCU2D add_2079_31 (.A0(resetn_c), .B0(n11558), .C0(quad_count[28]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[29]), 
          .D1(GND_net), .CIN(n25089), .COUT(n25090), .S0(n6366[28]), 
          .S1(n6366[29]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_31.INIT0 = 16'hd2d2;
    defparam add_2079_31.INIT1 = 16'hd2d2;
    defparam add_2079_31.INJECT1_0 = "NO";
    defparam add_2079_31.INJECT1_1 = "NO";
    CCU2D add_2079_29 (.A0(resetn_c), .B0(n11558), .C0(quad_count[26]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[27]), 
          .D1(GND_net), .CIN(n25088), .COUT(n25089), .S0(n6366[26]), 
          .S1(n6366[27]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_29.INIT0 = 16'hd2d2;
    defparam add_2079_29.INIT1 = 16'hd2d2;
    defparam add_2079_29.INJECT1_0 = "NO";
    defparam add_2079_29.INJECT1_1 = "NO";
    CCU2D add_2079_27 (.A0(resetn_c), .B0(n11558), .C0(quad_count[24]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[25]), 
          .D1(GND_net), .CIN(n25087), .COUT(n25088), .S0(n6366[24]), 
          .S1(n6366[25]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_27.INIT0 = 16'hd2d2;
    defparam add_2079_27.INIT1 = 16'hd2d2;
    defparam add_2079_27.INJECT1_0 = "NO";
    defparam add_2079_27.INJECT1_1 = "NO";
    CCU2D add_2079_25 (.A0(resetn_c), .B0(n11558), .C0(quad_count[22]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[23]), 
          .D1(GND_net), .CIN(n25086), .COUT(n25087), .S0(n6366[22]), 
          .S1(n6366[23]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_25.INIT0 = 16'hd2d2;
    defparam add_2079_25.INIT1 = 16'hd2d2;
    defparam add_2079_25.INJECT1_0 = "NO";
    defparam add_2079_25.INJECT1_1 = "NO";
    CCU2D add_2079_23 (.A0(resetn_c), .B0(n11558), .C0(quad_count[20]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[21]), 
          .D1(GND_net), .CIN(n25085), .COUT(n25086), .S0(n6366[20]), 
          .S1(n6366[21]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_23.INIT0 = 16'hd2d2;
    defparam add_2079_23.INIT1 = 16'hd2d2;
    defparam add_2079_23.INJECT1_0 = "NO";
    defparam add_2079_23.INJECT1_1 = "NO";
    CCU2D add_2079_21 (.A0(resetn_c), .B0(n11558), .C0(quad_count[18]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[19]), 
          .D1(GND_net), .CIN(n25084), .COUT(n25085), .S0(n6366[18]), 
          .S1(n6366[19]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_21.INIT0 = 16'hd2d2;
    defparam add_2079_21.INIT1 = 16'hd2d2;
    defparam add_2079_21.INJECT1_0 = "NO";
    defparam add_2079_21.INJECT1_1 = "NO";
    CCU2D add_2079_19 (.A0(resetn_c), .B0(n11558), .C0(quad_count[16]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[17]), 
          .D1(GND_net), .CIN(n25083), .COUT(n25084), .S0(n6366[16]), 
          .S1(n6366[17]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_19.INIT0 = 16'hd2d2;
    defparam add_2079_19.INIT1 = 16'hd2d2;
    defparam add_2079_19.INJECT1_0 = "NO";
    defparam add_2079_19.INJECT1_1 = "NO";
    CCU2D add_2079_17 (.A0(resetn_c), .B0(n11558), .C0(quad_count[14]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[15]), 
          .D1(GND_net), .CIN(n25082), .COUT(n25083), .S0(n6366[14]), 
          .S1(n6366[15]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_17.INIT0 = 16'hd2d2;
    defparam add_2079_17.INIT1 = 16'hd2d2;
    defparam add_2079_17.INJECT1_0 = "NO";
    defparam add_2079_17.INJECT1_1 = "NO";
    CCU2D add_2079_15 (.A0(resetn_c), .B0(n11558), .C0(quad_count[12]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[13]), 
          .D1(GND_net), .CIN(n25081), .COUT(n25082), .S0(n6366[12]), 
          .S1(n6366[13]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_15.INIT0 = 16'hd2d2;
    defparam add_2079_15.INIT1 = 16'hd2d2;
    defparam add_2079_15.INJECT1_0 = "NO";
    defparam add_2079_15.INJECT1_1 = "NO";
    CCU2D add_2079_13 (.A0(resetn_c), .B0(n11558), .C0(quad_count[10]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[11]), 
          .D1(GND_net), .CIN(n25080), .COUT(n25081), .S0(n6366[10]), 
          .S1(n6366[11]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_13.INIT0 = 16'hd2d2;
    defparam add_2079_13.INIT1 = 16'hd2d2;
    defparam add_2079_13.INJECT1_0 = "NO";
    defparam add_2079_13.INJECT1_1 = "NO";
    CCU2D add_2079_11 (.A0(resetn_c), .B0(n11558), .C0(quad_count[8]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[9]), 
          .D1(GND_net), .CIN(n25079), .COUT(n25080), .S0(n6366[8]), 
          .S1(n6366[9]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_11.INIT0 = 16'hd2d2;
    defparam add_2079_11.INIT1 = 16'hd2d2;
    defparam add_2079_11.INJECT1_0 = "NO";
    defparam add_2079_11.INJECT1_1 = "NO";
    CCU2D add_2079_9 (.A0(resetn_c), .B0(n11558), .C0(quad_count[6]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[7]), 
          .D1(GND_net), .CIN(n25078), .COUT(n25079), .S0(n6366[6]), 
          .S1(n6366[7]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_9.INIT0 = 16'hd2d2;
    defparam add_2079_9.INIT1 = 16'hd2d2;
    defparam add_2079_9.INJECT1_0 = "NO";
    defparam add_2079_9.INJECT1_1 = "NO";
    CCU2D add_2079_7 (.A0(resetn_c), .B0(n11558), .C0(quad_count[4]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[5]), 
          .D1(GND_net), .CIN(n25077), .COUT(n25078), .S0(n6366[4]), 
          .S1(n6366[5]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_7.INIT0 = 16'hd2d2;
    defparam add_2079_7.INIT1 = 16'hd2d2;
    defparam add_2079_7.INJECT1_0 = "NO";
    defparam add_2079_7.INJECT1_1 = "NO";
    CCU2D add_2079_5 (.A0(resetn_c), .B0(n11558), .C0(quad_count[2]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[3]), 
          .D1(GND_net), .CIN(n25076), .COUT(n25077), .S0(n6366[2]), 
          .S1(n6366[3]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_5.INIT0 = 16'hd2d2;
    defparam add_2079_5.INIT1 = 16'hd2d2;
    defparam add_2079_5.INJECT1_0 = "NO";
    defparam add_2079_5.INJECT1_1 = "NO";
    CCU2D add_2079_3 (.A0(resetn_c), .B0(n11558), .C0(quad_count[0]), 
          .D0(GND_net), .A1(resetn_c), .B1(n11558), .C1(quad_count[1]), 
          .D1(GND_net), .CIN(n25075), .COUT(n25076), .S0(n6366[0]), 
          .S1(n6366[1]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_3.INIT0 = 16'h2d2d;
    defparam add_2079_3.INIT1 = 16'hd2d2;
    defparam add_2079_3.INJECT1_0 = "NO";
    defparam add_2079_3.INJECT1_1 = "NO";
    CCU2D add_2079_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(resetn_c), .B1(n11558), .C1(GND_net), .D1(GND_net), .COUT(n25075));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_2079_1.INIT0 = 16'hF000;
    defparam add_2079_1.INIT1 = 16'hdddd;
    defparam add_2079_1.INJECT1_0 = "NO";
    defparam add_2079_1.INJECT1_1 = "NO";
    FD1S3AX quad_buffer_i31 (.D(quad_count[31]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i31.GSR = "DISABLED";
    FD1S3AX quad_buffer_i30 (.D(quad_count[30]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i30.GSR = "DISABLED";
    FD1S3AX quad_buffer_i29 (.D(quad_count[29]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i29.GSR = "DISABLED";
    FD1S3AX quad_buffer_i28 (.D(quad_count[28]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i28.GSR = "DISABLED";
    FD1S3AX quad_buffer_i27 (.D(quad_count[27]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i27.GSR = "DISABLED";
    FD1S3AX quad_buffer_i26 (.D(quad_count[26]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i26.GSR = "DISABLED";
    FD1S3AX quad_buffer_i25 (.D(quad_count[25]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i25.GSR = "DISABLED";
    FD1S3AX quad_buffer_i24 (.D(quad_count[24]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i24.GSR = "DISABLED";
    FD1S3AX quad_buffer_i23 (.D(quad_count[23]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i23.GSR = "DISABLED";
    FD1S3AX quad_buffer_i22 (.D(quad_count[22]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i22.GSR = "DISABLED";
    FD1S3AX quad_buffer_i21 (.D(quad_count[21]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i21.GSR = "DISABLED";
    FD1S3AX quad_buffer_i20 (.D(quad_count[20]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i20.GSR = "DISABLED";
    FD1S3AX quad_buffer_i19 (.D(quad_count[19]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i19.GSR = "DISABLED";
    FD1S3AX quad_buffer_i18 (.D(quad_count[18]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i18.GSR = "DISABLED";
    FD1S3AX quad_buffer_i17 (.D(quad_count[17]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i17.GSR = "DISABLED";
    FD1S3AX quad_buffer_i16 (.D(quad_count[16]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i16.GSR = "DISABLED";
    FD1S3AX quad_buffer_i15 (.D(quad_count[15]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i15.GSR = "DISABLED";
    FD1S3AX quad_buffer_i14 (.D(quad_count[14]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i14.GSR = "DISABLED";
    FD1S3AX quad_buffer_i13 (.D(quad_count[13]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i13.GSR = "DISABLED";
    FD1S3AX quad_buffer_i12 (.D(quad_count[12]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i12.GSR = "DISABLED";
    FD1S3AX quad_buffer_i11 (.D(quad_count[11]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i11.GSR = "DISABLED";
    FD1S3AX quad_buffer_i10 (.D(quad_count[10]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i10.GSR = "DISABLED";
    FD1S3AX quad_buffer_i9 (.D(quad_count[9]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i9.GSR = "DISABLED";
    FD1S3AX quad_buffer_i8 (.D(quad_count[8]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i8.GSR = "DISABLED";
    FD1S3AX quad_buffer_i7 (.D(quad_count[7]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i7.GSR = "DISABLED";
    FD1S3AX quad_buffer_i6 (.D(quad_count[6]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i6.GSR = "DISABLED";
    FD1S3AX quad_buffer_i5 (.D(quad_count[5]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i5.GSR = "DISABLED";
    FD1S3AX quad_buffer_i4 (.D(quad_count[4]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i4.GSR = "DISABLED";
    FD1S3AX quad_buffer_i3 (.D(quad_count[3]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i3.GSR = "DISABLED";
    FD1S3AX quad_buffer_i2 (.D(quad_count[2]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i2.GSR = "DISABLED";
    FD1S3AX quad_buffer_i1 (.D(quad_count[1]), .CK(\pin_intrpt[5] ), .Q(quad_buffer[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i1.GSR = "DISABLED";
    FD1S3AX AB_i1 (.D(sync[1]), .CK(clk_1MHz), .Q(AB[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam AB_i1.GSR = "DISABLED";
    FD1S3AX sync_i1 (.D(\quad_a[1] ), .CK(clk_1MHz), .Q(sync[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam sync_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_1313[31] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i31 (.D(\spi_data_out_r_39__N_1313[30] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i30 (.D(\spi_data_out_r_39__N_1313[29] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i29 (.D(\spi_data_out_r_39__N_1313[28] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i28 (.D(\spi_data_out_r_39__N_1313[27] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i27 (.D(\spi_data_out_r_39__N_1313[26] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i26 (.D(\spi_data_out_r_39__N_1313[25] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i25 (.D(\spi_data_out_r_39__N_1313[24] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i24 (.D(\spi_data_out_r_39__N_1313[23] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i23 (.D(\spi_data_out_r_39__N_1313[22] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i22 (.D(\spi_data_out_r_39__N_1313[21] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i21 (.D(\spi_data_out_r_39__N_1313[20] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i20 (.D(\spi_data_out_r_39__N_1313[19] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i19 (.D(\spi_data_out_r_39__N_1313[18] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i18 (.D(\spi_data_out_r_39__N_1313[17] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i17 (.D(\spi_data_out_r_39__N_1313[16] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i16 (.D(\spi_data_out_r_39__N_1313[15] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_1313[14] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_1313[13] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_1313[12] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_1313[11] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_1313[10] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_1313[9] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_1313[8] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_1313[7] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_1313[6] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_1313[5] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_1313[4] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_1313[3] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_1313[2] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_1313[1] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_1168[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i31 (.D(n25837), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i31.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i30 (.D(n25835), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i30.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i29 (.D(n25857), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i29.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i28 (.D(n25855), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i28.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i27 (.D(n25877), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i27.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i26 (.D(n25875), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i26.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i25 (.D(n25897), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i25.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i24 (.D(n25895), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i24.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i23 (.D(n25917), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i23.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i22 (.D(n25915), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i22.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i21 (.D(n25937), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i21.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i20 (.D(n25935), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i20.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i19 (.D(n25957), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i19.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i18 (.D(n25955), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i18.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i17 (.D(n25977), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i17.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i16 (.D(n25975), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i16.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i15 (.D(n25997), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i15.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i14 (.D(n25995), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i14.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i13 (.D(n26017), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i13.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i12 (.D(n26015), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i12.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i11 (.D(n26037), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i11.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i10 (.D(n26035), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i10.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i9 (.D(n26065), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i9.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i8 (.D(n26063), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i8.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i7 (.D(n26091), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i7.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i6 (.D(n26089), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i6.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i5 (.D(n26111), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i5.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i4 (.D(n26109), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i4.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i3 (.D(n26139), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i3.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i2 (.D(n26137), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i1 (.D(n26167), .SP(clk_1MHz_enable_309), .CK(clk_1MHz), 
            .Q(quad_count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i1.GSR = "DISABLED";
    FD1P3IX quad_homing__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_286), .CD(n29239), 
            .CK(clk), .Q(\quad_homing[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam quad_homing__i1.GSR = "DISABLED";
    FD1P3IX quad_set__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i1.GSR = "DISABLED";
    FD1P3IX quad_set__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i2.GSR = "DISABLED";
    FD1P3IX quad_set__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i3.GSR = "DISABLED";
    FD1P3IX quad_set__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i4.GSR = "DISABLED";
    FD1P3IX quad_set__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i5.GSR = "DISABLED";
    FD1P3IX quad_set__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i6.GSR = "DISABLED";
    FD1P3IX quad_set__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i7.GSR = "DISABLED";
    FD1P3IX quad_set__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i8.GSR = "DISABLED";
    FD1P3IX quad_set__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i9.GSR = "DISABLED";
    FD1P3IX quad_set__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i10.GSR = "DISABLED";
    FD1P3IX quad_set__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i11.GSR = "DISABLED";
    FD1P3IX quad_set__i12 (.D(\spi_data_r[12] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i12.GSR = "DISABLED";
    FD1P3IX quad_set__i13 (.D(\spi_data_r[13] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i13.GSR = "DISABLED";
    FD1P3IX quad_set__i14 (.D(\spi_data_r[14] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i14.GSR = "DISABLED";
    FD1P3IX quad_set__i15 (.D(\spi_data_r[15] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i15.GSR = "DISABLED";
    FD1P3IX quad_set__i16 (.D(\spi_data_r[16] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i16.GSR = "DISABLED";
    FD1P3IX quad_set__i17 (.D(\spi_data_r[17] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i17.GSR = "DISABLED";
    FD1P3IX quad_set__i18 (.D(\spi_data_r[18] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i18.GSR = "DISABLED";
    FD1P3IX quad_set__i19 (.D(\spi_data_r[19] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i19.GSR = "DISABLED";
    FD1P3IX quad_set__i20 (.D(\spi_data_r[20] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i20.GSR = "DISABLED";
    FD1P3IX quad_set__i21 (.D(\spi_data_r[21] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i21.GSR = "DISABLED";
    FD1P3IX quad_set__i22 (.D(\spi_data_r[22] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i22.GSR = "DISABLED";
    FD1P3IX quad_set__i23 (.D(\spi_data_r[23] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i23.GSR = "DISABLED";
    FD1P3IX quad_set__i24 (.D(\spi_data_r[24] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i24.GSR = "DISABLED";
    FD1P3IX quad_set__i25 (.D(\spi_data_r[25] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i25.GSR = "DISABLED";
    FD1P3IX quad_set__i26 (.D(\spi_data_r[26] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i26.GSR = "DISABLED";
    FD1P3IX quad_set__i27 (.D(\spi_data_r[27] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i27.GSR = "DISABLED";
    FD1P3IX quad_set__i28 (.D(\spi_data_r[28] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i28.GSR = "DISABLED";
    FD1P3IX quad_set__i29 (.D(\spi_data_r[29] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i29.GSR = "DISABLED";
    FD1P3IX quad_set__i30 (.D(\spi_data_r[30] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i30.GSR = "DISABLED";
    FD1P3IX quad_set__i31 (.D(\spi_data_r[31] ), .SP(clk_enable_467), .CD(n29239), 
            .CK(clk), .Q(quad_set[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i31.GSR = "DISABLED";
    LUT4 i31_4_lut (.A(n6366[31]), .B(quad_set[31]), .C(n3), .D(n27061), 
         .Z(n25837)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut.init = 16'hcac0;
    LUT4 i31_4_lut_adj_808 (.A(n6366[30]), .B(quad_set[30]), .C(n3), .D(n27061), 
         .Z(n25835)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_808.init = 16'hcac0;
    LUT4 i31_4_lut_adj_809 (.A(n6366[29]), .B(quad_set[29]), .C(n3), .D(n27061), 
         .Z(n25857)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_809.init = 16'hcac0;
    LUT4 i31_4_lut_adj_810 (.A(n6366[28]), .B(quad_set[28]), .C(n3), .D(n27061), 
         .Z(n25855)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_810.init = 16'hcac0;
    LUT4 i31_4_lut_adj_811 (.A(n6366[27]), .B(quad_set[27]), .C(n3), .D(n27061), 
         .Z(n25877)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_811.init = 16'hcac0;
    LUT4 i31_4_lut_adj_812 (.A(n6366[26]), .B(quad_set[26]), .C(n3), .D(n27061), 
         .Z(n25875)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_812.init = 16'hcac0;
    FD1P3IX quad_set_valid_404 (.D(n29084), .SP(clk_enable_502), .CD(n29239), 
            .CK(clk), .Q(quad_set_valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set_valid_404.GSR = "DISABLED";
    LUT4 i31_4_lut_adj_813 (.A(n6366[25]), .B(quad_set[25]), .C(n3), .D(n27061), 
         .Z(n25897)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_813.init = 16'hcac0;
    LUT4 i31_4_lut_adj_814 (.A(n6366[24]), .B(quad_set[24]), .C(n3), .D(n27061), 
         .Z(n25895)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_814.init = 16'hcac0;
    LUT4 i31_4_lut_adj_815 (.A(n6366[23]), .B(quad_set[23]), .C(n3), .D(n27061), 
         .Z(n25917)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_815.init = 16'hcac0;
    LUT4 i31_4_lut_adj_816 (.A(n6366[22]), .B(quad_set[22]), .C(n3), .D(n27061), 
         .Z(n25915)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_816.init = 16'hcac0;
    LUT4 i31_4_lut_adj_817 (.A(n6366[21]), .B(quad_set[21]), .C(n3), .D(n27061), 
         .Z(n25937)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_817.init = 16'hcac0;
    LUT4 i31_4_lut_adj_818 (.A(n6366[20]), .B(quad_set[20]), .C(n3), .D(n27061), 
         .Z(n25935)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_818.init = 16'hcac0;
    LUT4 i31_4_lut_adj_819 (.A(n6366[19]), .B(quad_set[19]), .C(n3), .D(n27061), 
         .Z(n25957)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_819.init = 16'hcac0;
    LUT4 i31_4_lut_adj_820 (.A(n6366[18]), .B(quad_set[18]), .C(n3), .D(n27061), 
         .Z(n25955)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_820.init = 16'hcac0;
    LUT4 i31_4_lut_adj_821 (.A(n6366[17]), .B(quad_set[17]), .C(n3), .D(n27061), 
         .Z(n25977)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_821.init = 16'hcac0;
    LUT4 i31_4_lut_adj_822 (.A(n6366[16]), .B(quad_set[16]), .C(n3), .D(n27061), 
         .Z(n25975)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_822.init = 16'hcac0;
    LUT4 i31_4_lut_adj_823 (.A(n6366[15]), .B(quad_set[15]), .C(n3), .D(n27061), 
         .Z(n25997)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_823.init = 16'hcac0;
    LUT4 i31_4_lut_adj_824 (.A(n6366[14]), .B(quad_set[14]), .C(n3), .D(n27061), 
         .Z(n25995)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_824.init = 16'hcac0;
    LUT4 i31_4_lut_adj_825 (.A(n6366[13]), .B(quad_set[13]), .C(n3), .D(n27061), 
         .Z(n26017)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_825.init = 16'hcac0;
    LUT4 i31_4_lut_adj_826 (.A(n6366[12]), .B(quad_set[12]), .C(n3), .D(n27061), 
         .Z(n26015)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_826.init = 16'hcac0;
    LUT4 i31_4_lut_adj_827 (.A(n6366[11]), .B(quad_set[11]), .C(n3), .D(n27061), 
         .Z(n26037)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_827.init = 16'hcac0;
    LUT4 i31_4_lut_adj_828 (.A(n6366[10]), .B(quad_set[10]), .C(n3), .D(n27061), 
         .Z(n26035)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_828.init = 16'hcac0;
    LUT4 i31_4_lut_adj_829 (.A(n6366[9]), .B(quad_set[9]), .C(n3), .D(n27061), 
         .Z(n26065)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_829.init = 16'hcac0;
    LUT4 i31_4_lut_adj_830 (.A(n6366[8]), .B(quad_set[8]), .C(n3), .D(n27061), 
         .Z(n26063)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_830.init = 16'hcac0;
    LUT4 i31_4_lut_adj_831 (.A(n6366[7]), .B(quad_set[7]), .C(n3), .D(n27061), 
         .Z(n26091)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_831.init = 16'hcac0;
    LUT4 i31_4_lut_adj_832 (.A(n6366[6]), .B(quad_set[6]), .C(n3), .D(n27061), 
         .Z(n26089)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_832.init = 16'hcac0;
    LUT4 i31_4_lut_adj_833 (.A(n6366[5]), .B(quad_set[5]), .C(n3), .D(n27061), 
         .Z(n26111)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_833.init = 16'hcac0;
    LUT4 i31_4_lut_adj_834 (.A(n6366[4]), .B(quad_set[4]), .C(n3), .D(n27061), 
         .Z(n26109)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_834.init = 16'hcac0;
    LUT4 i31_4_lut_adj_835 (.A(n6366[3]), .B(quad_set[3]), .C(n3), .D(n27061), 
         .Z(n26139)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_835.init = 16'hcac0;
    LUT4 i31_4_lut_adj_836 (.A(n6366[2]), .B(quad_set[2]), .C(n3), .D(n27061), 
         .Z(n26137)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_836.init = 16'hcac0;
    LUT4 i31_4_lut_adj_837 (.A(n6366[1]), .B(quad_set[1]), .C(n3), .D(n27061), 
         .Z(n26167)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_837.init = 16'hcac0;
    LUT4 i22938_4_lut (.A(quad_set_valid), .B(resetn_c), .C(n26753), .D(n12716), 
         .Z(clk_1MHz_enable_309)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i22938_4_lut.init = 16'hffbf;
    LUT4 i31_4_lut_adj_838 (.A(n6366[0]), .B(quad_set[0]), .C(n3), .D(n27061), 
         .Z(n26141)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i31_4_lut_adj_838.init = 16'hcac0;
    LUT4 i2_4_lut (.A(n26963), .B(quad_set_valid), .C(n4), .D(resetn_c), 
         .Z(n3)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'h8000;
    LUT4 i1_3_lut (.A(resetn_c), .B(n12716), .C(n4), .Z(n27061)) /* synthesis lut_function=(!((B (C))+!A)) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i1_3_lut.init = 16'h2a2a;
    LUT4 i1_4_lut (.A(n1521[1]), .B(n12), .C(n1521[2]), .D(n1521[3]), 
         .Z(n4)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i1_4_lut.init = 16'h33c9;
    LUT4 i15_2_lut (.A(AB[1]), .B(AB[0]), .Z(n12)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(155[16] 158[10])
    defparam i15_2_lut.init = 16'h6666;
    LUT4 i22466_2_lut (.A(quad_homing[0]), .B(pin_io_out_14), .Z(n27636)) /* synthesis lut_function=(A (B)) */ ;
    defparam i22466_2_lut.init = 16'h8888;
    LUT4 i1_2_lut (.A(n1521[1]), .B(n1521[2]), .Z(n8)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_adj_839 (.A(n1521[0]), .B(n1521[3]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam i1_2_lut_adj_839.init = 16'heeee;
    LUT4 n8_bdd_4_lut (.A(n8), .B(n1521[0]), .C(AB[1]), .D(AB[0]), .Z(n28864)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D)))) */ ;
    defparam n8_bdd_4_lut.init = 16'hc00e;
    
endmodule
//
// Verilog Description of module \stepper(DEV_ID=6,UART_ADDRESS_WIDTH=4) 
//

module \stepper(DEV_ID=6,UART_ADDRESS_WIDTH=4)  (\spi_data_out_r[26] , \spi_data_out_r_39__N_1168[26] , 
            spi_data_out_r_39__N_1208, mode_adj_181, clk, clk_enable_288, 
            n29239, n29762, \spi_data_out_r_39__N_1636[15] , spi_data_out_r_39__N_1676, 
            \spi_data_out_r_39__N_4835[26] , spi_data_out_r_39__N_4875, 
            \spi_data_out_r_39__N_5513[26] , spi_data_out_r_39__N_5553, 
            \spi_data_out_r_39__N_4496[26] , spi_data_out_r_39__N_4536, 
            \spi_data_out_r_39__N_3818[26] , spi_data_out_r_39__N_3858, 
            \spi_data_out_r_39__N_2104[26] , \spi_data_out_r_39__N_1870[26] , 
            spi_data_out_r_39__N_2144, spi_data_out_r_39__N_1910, \spi_data_out_r_39__N_1402[26] , 
            spi_data_out_r_39__N_1442, \spi_data_out_r_39__N_2338[26] , 
            \spi_data_out_r_39__N_5174[26] , spi_data_out_r_39__N_2378, 
            spi_data_out_r_39__N_5214, \spi_data_out_r_39__N_1636[26] , 
            \spi_data_out_r_39__N_934[26] , spi_data_out_r_39__N_974, spi_data_out_r_39__N_5892, 
            \spi_data_out_r_39__N_4157[26] , spi_data_out_r_39__N_4197, 
            pin_io_out_68, \quad_a[6] , n28811, \spi_data_out_r[27] , 
            pin_io_out_69, \quad_b[6] , \spi_data_out_r_39__N_1168[27] , 
            \spi_data_out_r_39__N_4835[27] , \spi_data_out_r_39__N_5513[27] , 
            \spi_data_out_r_39__N_4835[21] , \spi_data_out_r_39__N_4496[27] , 
            \spi_data_out_r_39__N_3818[27] , \spi_data_out_r_39__N_2104[27] , 
            \spi_data_out_r_39__N_1870[27] , \spi_data_out_r_39__N_1402[27] , 
            \spi_data_out_r_39__N_2338[27] , \spi_data_out_r_39__N_5174[27] , 
            \spi_data_out_r_39__N_1636[27] , \spi_data_out_r_39__N_934[27] , 
            \spi_data_out_r_39__N_4157[27] , \spi_data_out_r[28] , \spi_data_out_r_39__N_1168[28] , 
            \SLO_buf[0] , \spi_data_out_r_39__N_5852[0] , \spi_data_out_r_39__N_6114[0] , 
            \spi_data_out_r_39__N_4835[28] , clk_1MHz, clk_1MHz_enable_367, 
            \spi_data_out_r_39__N_5513[28] , \spi_data_out_r_39__N_934[15] , 
            \spi_data_out_r_39__N_4157[15] , \spi_data_out_r_39__N_4496[28] , 
            \spi_data_out_r_39__N_3818[28] , \spi_data_out_r_39__N_2104[28] , 
            \spi_data_out_r_39__N_1870[28] , \spi_data_out_r_39__N_1402[28] , 
            \spi_data_out_r_39__N_2338[28] , \spi_data_out_r_39__N_5174[28] , 
            \spi_data_out_r_39__N_1636[21] , \spi_data_out_r_39__N_934[21] , 
            \spi_data_out_r_39__N_4157[21] , \spi_data_out_r_39__N_1636[28] , 
            \spi_data_out_r[22] , \spi_data_out_r_39__N_1168[22] , \spi_data_out_r_39__N_4835[22] , 
            \spi_data_out_r_39__N_5513[22] , \spi_data_out_r_39__N_934[28] , 
            \spi_data_out_r_39__N_4157[28] , \spi_data_out_r[29] , \spi_data_out_r_39__N_4496[22] , 
            \spi_data_out_r_39__N_1168[29] , \spi_data_out_r_39__N_4835[29] , 
            \spi_data_out_r_39__N_5513[29] , \spi_data_out_r_39__N_4496[29] , 
            \spi_data_out_r_39__N_3818[29] , \spi_data_out_r_39__N_3818[22] , 
            \spi_data_out_r_39__N_2104[29] , \spi_data_out_r_39__N_1870[29] , 
            \spi_data_out_r_39__N_2104[22] , \spi_data_out_r_39__N_1870[22] , 
            \spi_data_out_r_39__N_1402[22] , \spi_data_out_r_39__N_1402[29] , 
            \spi_data_out_r_39__N_2338[29] , \spi_data_out_r_39__N_5174[29] , 
            \spi_data_out_r_39__N_1636[29] , \spi_data_out_r_39__N_2338[22] , 
            \spi_data_out_r_39__N_5174[22] , \spi_data_out_r_39__N_934[29] , 
            n29087, \spi_data_out_r_39__N_4157[29] , \spi_data_out_r_39__N_1636[22] , 
            \spi_data_out_r[30] , \spi_data_out_r_39__N_1168[30] , \spi_data_out_r_39__N_934[22] , 
            \spi_data_out_r_39__N_4835[30] , \spi_data_out_r_39__N_5513[30] , 
            \spi_data_out_r_39__N_4157[22] , \spi_data_out_r_39__N_4496[30] , 
            \spi_data_out_r[23] , \spi_data_out_r_39__N_3818[30] , digital_output_r, 
            clk_enable_198, \spi_data_r[0] , \spi_data_out_r_39__N_1168[23] , 
            \spi_data_out_r_39__N_2104[30] , \spi_data_out_r_39__N_1870[30] , 
            \spi_data_out_r_39__N_1402[30] , \spi_data_out_r_39__N_2338[30] , 
            \spi_data_out_r_39__N_5174[30] , \spi_data_out_r_39__N_1636[30] , 
            \spi_data_out_r_39__N_934[30] , \spi_data_out_r_39__N_4157[30] , 
            \spi_data_out_r[31] , \spi_data_out_r_39__N_4835[23] , \spi_data_out_r_39__N_1168[31] , 
            \spi_data_out_r_39__N_5513[23] , \spi_data_out_r[16] , \spi_data_out_r_39__N_1168[16] , 
            \spi_data_out_r_39__N_4496[23] , \spi_data_out_r_39__N_4835[31] , 
            \spi_data_out_r_39__N_3818[23] , \spi_data_out_r_39__N_5513[31] , 
            \spi_data_out_r_39__N_4496[31] , n19401, resetn_c, \spi_data_out_r_39__N_3818[31] , 
            \spi_data_out_r_39__N_2104[31] , \spi_data_out_r_39__N_1870[31] , 
            \spi_data_out_r_39__N_1402[31] , \spi_data_out_r_39__N_2338[31] , 
            \spi_data_out_r_39__N_5174[31] , \spi_data_out_r_39__N_1636[31] , 
            \spi_data_out_r_39__N_934[31] , \spi_data_out_r_39__N_4157[31] , 
            \spi_data_out_r_39__N_4835[32] , \spi_data_out_r[32] , \spi_data_out_r_39__N_3818[32] , 
            \spi_data_out_r_39__N_5174[32] , \spi_data_out_r_39__N_4496[32] , 
            \spi_data_out_r_39__N_4157[32] , \spi_data_out_r_39__N_5513[32] , 
            \spi_data_out_r_39__N_4835[33] , \spi_data_out_r[33] , \spi_data_out_r_39__N_3818[33] , 
            \spi_data_out_r_39__N_5174[33] , \spi_data_out_r_39__N_4496[33] , 
            \spi_data_out_r_39__N_4157[33] , \spi_data_out_r_39__N_5513[33] , 
            \spi_data_out_r_39__N_4835[34] , \spi_data_out_r[34] , \spi_data_out_r_39__N_3818[34] , 
            \spi_data_out_r_39__N_5174[34] , \spi_data_out_r_39__N_4496[34] , 
            \spi_data_out_r_39__N_4157[34] , \spi_data_out_r_39__N_2104[23] , 
            \spi_data_out_r_39__N_1870[23] , \spi_data_out_r_39__N_5513[34] , 
            \spi_data_out_r_39__N_4835[35] , \spi_data_out_r[35] , \spi_data_out_r_39__N_3818[35] , 
            \spi_data_out_r_39__N_5174[35] , \spi_data_out_r_39__N_4496[35] , 
            \spi_data_out_r_39__N_4157[35] , \spi_data_out_r_39__N_5513[35] , 
            \spi_data_out_r_39__N_4835[36] , \spi_data_out_r[36] , \spi_data_out_r_39__N_3818[36] , 
            \spi_data_out_r_39__N_5174[36] , \spi_data_out_r_39__N_4496[36] , 
            \spi_data_out_r_39__N_4157[36] , \spi_data_out_r_39__N_5513[36] , 
            \spi_data_out_r_39__N_4835[37] , \spi_data_out_r[37] , \spi_data_out_r_39__N_1402[23] , 
            \spi_data_out_r_39__N_3818[37] , \spi_data_out_r_39__N_5174[37] , 
            \spi_data_out_r_39__N_4496[37] , \spi_data_out_r_39__N_4157[37] , 
            \spi_data_out_r_39__N_2338[23] , \spi_data_out_r_39__N_5174[23] , 
            \spi_data_out_r_39__N_5513[37] , \spi_data_out_r_39__N_4835[38] , 
            \spi_data_out_r[38] , \spi_data_out_r_39__N_3818[38] , \spi_data_out_r_39__N_1636[23] , 
            \spi_data_out_r_39__N_5174[38] , \spi_data_out_r_39__N_4496[38] , 
            \spi_data_out_r_39__N_4157[38] , \spi_data_out_r_39__N_934[23] , 
            \spi_data_out_r_39__N_4157[23] , \spi_data_out_r_39__N_5513[38] , 
            \spi_data_out_r_39__N_4835[39] , \spi_data_out_r[39] , \spi_data_out_r_39__N_3818[39] , 
            \spi_data_out_r_39__N_5174[39] , \spi_data_out_r_39__N_4496[39] , 
            \spi_data_out_r_39__N_4157[39] , \spi_data_out_r_39__N_5513[39] , 
            \spi_data_out_r[24] , \spi_data_out_r_39__N_1168[24] , \spi_data_out_r_39__N_4835[24] , 
            \spi_data_out_r_39__N_5513[24] , \spi_data_out_r_39__N_4496[24] , 
            n29267, mode, n29191, n29153, \spi_data_out_r_39__N_3818[24] , 
            n29195, \spi_data_out_r_39__N_2104[24] , \spi_data_out_r_39__N_1870[24] , 
            n29293, \cs_decoded[12] , n8652, n1, n8651, n1_adj_171, 
            \spi_data_out_r_39__N_5513[21] , \spi_data_out_r_39__N_1402[24] , 
            \spi_data_out_r_39__N_2338[24] , \spi_data_out_r_39__N_5174[24] , 
            \spi_data_out_r_39__N_1636[24] , \spi_data_out_r_39__N_934[24] , 
            \spi_data_out_r_39__N_4157[24] , \spi_data_out_r[25] , \spi_data_out_r_39__N_1168[25] , 
            \spi_data_out_r_39__N_4835[25] , \spi_data_out_r_39__N_5513[25] , 
            \spi_data_out_r_39__N_4496[25] , \spi_data_out_r_39__N_3818[25] , 
            \spi_data_out_r_39__N_2104[25] , \spi_data_out_r_39__N_1870[25] , 
            \spi_data_out_r_39__N_1402[25] , \spi_data_out_r_39__N_2338[25] , 
            \spi_data_out_r_39__N_5174[25] , GND_net, \spi_data_out_r_39__N_1636[25] , 
            \spi_data_out_r_39__N_934[25] , \spi_data_out_r_39__N_4157[25] , 
            \spi_data_r[2] , \spi_data_r[1] , \spi_data_out_r_39__N_4835[16] , 
            \spi_data_out_r_39__N_2856[2] , clear_intrpt, n13, \spi_data_out_r_39__N_1402[2] , 
            n4, \SLO_buf[1] , \SLO_buf[2] , \SLO_buf[3] , \SLO_buf[4] , 
            \SLO_buf[5] , \SLO_buf[6] , \SLO_buf[7] , \SLO_buf[8] , 
            \SLO_buf[9] , \SLO_buf[10] , \SLO_buf[11] , \SLO_buf[12] , 
            \SLO_buf[13] , \SLO_buf[14] , \SLO_buf[15] , \SLO_buf[16] , 
            \SLO_buf[17] , \SLO_buf[18] , \SLO_buf[19] , \SLO_buf[20] , 
            \SLO_buf[21] , \SLO_buf[22] , \SLO_buf[23] , \SLO_buf[24] , 
            \SLO_buf[25] , \SLO_buf[26] , \SLO_buf[27] , \SLO_buf[28] , 
            \SLO_buf[29] , \spi_data_out_r_39__N_5513[16] , \spi_data_out_r_39__N_6114[1] , 
            \spi_data_out_r_39__N_5852[2] , \spi_data_out_r_39__N_6114[2] , 
            \spi_data_out_r_39__N_6114[3] , \spi_data_out_r_39__N_6114[4] , 
            \spi_data_out_r_39__N_6114[5] , \spi_data_out_r_39__N_6114[6] , 
            \spi_data_out_r_39__N_6114[7] , \spi_data_out_r_39__N_6114[8] , 
            \spi_data_out_r_39__N_6114[9] , \spi_data_out_r_39__N_6114[10] , 
            \spi_data_out_r_39__N_6114[11] , \spi_data_out_r_39__N_6114[12] , 
            \spi_data_out_r_39__N_6114[13] , \spi_data_out_r_39__N_6114[14] , 
            \spi_data_out_r_39__N_6114[15] , n29076, \spi_data_out_r_39__N_6114[32] , 
            \spi_data_out_r_39__N_6114[33] , \spi_data_out_r_39__N_6114[34] , 
            \spi_data_out_r_39__N_6114[35] , \spi_data_out_r_39__N_4496[16] , 
            \spi_data_out_r_39__N_2338[2] , n8, \spi_data_out_r_39__N_2998[2] , 
            clear_intrpt_adj_172, n15, \spi_data_out_r_39__N_2714[2] , 
            clear_intrpt_adj_173, n11, \spi_data_out_r_39__N_4835[2] , 
            n19, \spi_data_out_r_39__N_3818[16] , \spi_data_out_r_39__N_4157[0] , 
            n17, \spi_data_out_r_39__N_1168[0] , n3, \spi_data_out_r_39__N_5174[0] , 
            n20, \spi_data_out_r_39__N_2998[0] , n15_adj_174, \spi_data_out_r_39__N_934[0] , 
            n2, \spi_data_out_r_39__N_5513[0] , n21, \spi_data_out_r_39__N_1402[0] , 
            n4_adj_175, \spi_data_out_r_39__N_2714[0] , n11_adj_176, \spi_data_out_r[1] , 
            \spi_data_out_r_39__N_2643[1] , \spi_data_out_r_39__N_2856[1] , 
            clear_intrpt_adj_177, \spi_data_out_r_39__N_934[1] , \spi_data_out_r_39__N_4157[1] , 
            \spi_data_out_r_39__N_1168[1] , \spi_data_out_r_39__N_2927[1] , 
            \spi_data_out_r_39__N_2785[1] , clear_intrpt_adj_178, clear_intrpt_adj_179, 
            \spi_data_out_r_39__N_1402[1] , \spi_data_out_r_39__N_5174[1] , 
            \spi_data_out_r_39__N_3818[1] , \spi_data_out_r_39__N_2338[1] , 
            \spi_data_out_r_39__N_4496[21] , \spi_data_out_r_39__N_4496[1] , 
            \spi_data_out_r_39__N_1870[1] , \spi_data_out_r_39__N_2998[1] , 
            \spi_data_out_r_39__N_2104[1] , \spi_data_out_r_39__N_2572[1] , 
            clear_intrpt_adj_180, \spi_data_out_r_39__N_4835[1] , \spi_data_out_r_39__N_5513[1] , 
            \spi_data_out_r_39__N_1636[1] , \spi_data_out_r_39__N_2714[1] , 
            \spi_data_out_r[3] , \spi_data_out_r_39__N_1168[3] , \spi_data_out_r_39__N_4835[3] , 
            \spi_data_out_r_39__N_5513[3] , \spi_data_out_r_39__N_4496[3] , 
            \spi_data_out_r_39__N_3818[3] , \spi_data_out_r_39__N_2104[3] , 
            \spi_data_out_r_39__N_1870[3] , \spi_data_out_r_39__N_1402[3] , 
            \spi_data_out_r_39__N_2338[3] , \spi_data_out_r_39__N_5174[3] , 
            \spi_data_out_r_39__N_1636[3] , \spi_data_out_r_39__N_934[3] , 
            \spi_data_out_r_39__N_4157[3] , \spi_data_out_r[4] , \spi_data_out_r_39__N_1168[4] , 
            \spi_data_out_r_39__N_4835[4] , \spi_data_out_r_39__N_5513[4] , 
            \spi_data_out_r_39__N_4496[4] , \spi_data_out_r_39__N_2104[16] , 
            \spi_data_out_r_39__N_1870[16] , \spi_data_out_r_39__N_3818[4] , 
            \spi_data_out_r_39__N_2104[4] , \spi_data_out_r_39__N_1870[4] , 
            \spi_data_out_r_39__N_1402[16] , \spi_data_out_r_39__N_1402[4] , 
            \spi_data_out_r_39__N_2338[4] , \spi_data_out_r_39__N_5174[4] , 
            \spi_data_out_r_39__N_1636[4] , \spi_data_out_r_39__N_934[4] , 
            \spi_data_out_r_39__N_4157[4] , \spi_data_out_r[5] , \spi_data_out_r_39__N_1168[5] , 
            \spi_data_out_r_39__N_4835[5] , \spi_data_out_r_39__N_5513[5] , 
            \spi_data_out_r_39__N_4496[5] , \spi_data_out_r_39__N_3818[5] , 
            \spi_data_out_r_39__N_2104[5] , \spi_data_out_r_39__N_1870[5] , 
            \spi_data_out_r_39__N_1402[5] , \spi_data_out_r_39__N_2338[5] , 
            \spi_data_out_r_39__N_5174[5] , \spi_data_out_r_39__N_1636[5] , 
            \spi_data_out_r_39__N_934[5] , \spi_data_out_r_39__N_4157[5] , 
            \spi_data_out_r[6] , \spi_data_out_r_39__N_1168[6] , \spi_data_out_r_39__N_4835[6] , 
            \spi_data_out_r_39__N_5513[6] , \spi_data_out_r_39__N_4496[6] , 
            \spi_data_out_r_39__N_3818[6] , \spi_data_out_r_39__N_2104[6] , 
            \spi_data_out_r_39__N_1870[6] , \spi_data_out_r_39__N_1402[6] , 
            \spi_data_out_r_39__N_2338[6] , \spi_data_out_r_39__N_5174[6] , 
            \spi_data_out_r_39__N_1636[6] , \spi_data_out_r_39__N_934[6] , 
            \spi_data_out_r_39__N_4157[6] , \spi_data_out_r[7] , \spi_data_out_r_39__N_1168[7] , 
            \spi_data_out_r_39__N_4835[7] , \spi_data_out_r_39__N_5513[7] , 
            \spi_data_out_r_39__N_4496[7] , \spi_data_out_r_39__N_3818[7] , 
            \spi_data_out_r_39__N_2104[7] , \spi_data_out_r_39__N_1870[7] , 
            \spi_data_out_r_39__N_1402[7] , \spi_data_out_r_39__N_2338[7] , 
            \spi_data_out_r_39__N_5174[7] , \spi_data_out_r_39__N_1636[7] , 
            \spi_data_out_r_39__N_934[7] , \spi_data_out_r_39__N_4157[7] , 
            \spi_data_out_r[8] , \spi_data_out_r_39__N_1168[8] , \spi_data_out_r_39__N_4835[8] , 
            \spi_data_out_r_39__N_5513[8] , \spi_data_out_r_39__N_4496[8] , 
            \spi_data_out_r_39__N_3818[8] , \spi_data_out_r_39__N_2104[8] , 
            \spi_data_out_r_39__N_1870[8] , \spi_data_out_r_39__N_1402[8] , 
            \spi_data_out_r_39__N_2338[8] , \spi_data_out_r_39__N_5174[8] , 
            \spi_data_out_r_39__N_1636[8] , \spi_data_out_r_39__N_934[8] , 
            \spi_data_out_r_39__N_4157[8] , \spi_data_out_r[9] , \spi_data_out_r_39__N_1168[9] , 
            \spi_data_out_r_39__N_4835[9] , \spi_data_out_r_39__N_5513[9] , 
            \spi_data_out_r_39__N_4496[9] , \spi_data_out_r_39__N_3818[9] , 
            \spi_data_out_r_39__N_2104[9] , \spi_data_out_r_39__N_1870[9] , 
            \spi_data_out_r_39__N_1402[9] , \spi_data_out_r_39__N_2338[9] , 
            \spi_data_out_r_39__N_5174[9] , \spi_data_out_r_39__N_1636[9] , 
            \spi_data_out_r_39__N_2338[16] , \spi_data_out_r_39__N_5174[16] , 
            \spi_data_out_r_39__N_934[9] , \spi_data_out_r_39__N_4157[9] , 
            \spi_data_out_r[10] , \spi_data_out_r_39__N_1168[10] , \spi_data_out_r_39__N_4835[10] , 
            \spi_data_out_r_39__N_5513[10] , \spi_data_out_r_39__N_4496[10] , 
            \spi_data_out_r_39__N_3818[10] , \spi_data_out_r_39__N_2104[10] , 
            \spi_data_out_r_39__N_1870[10] , \spi_data_out_r_39__N_1402[10] , 
            \spi_data_out_r_39__N_2338[10] , \spi_data_out_r_39__N_5174[10] , 
            \spi_data_out_r_39__N_1636[10] , \spi_data_out_r_39__N_934[10] , 
            \spi_data_out_r_39__N_4157[10] , \spi_data_out_r[11] , \spi_data_out_r_39__N_1168[11] , 
            \spi_data_out_r_39__N_4835[11] , \spi_data_out_r_39__N_5513[11] , 
            \spi_data_out_r_39__N_4496[11] , \spi_data_out_r_39__N_3818[11] , 
            \spi_data_out_r_39__N_2104[11] , \spi_data_out_r_39__N_1870[11] , 
            \spi_data_out_r_39__N_1402[11] , \spi_data_out_r_39__N_2338[11] , 
            \spi_data_out_r_39__N_5174[11] , \spi_data_out_r_39__N_1636[11] , 
            \spi_data_out_r_39__N_934[11] , \spi_data_out_r_39__N_4157[11] , 
            \spi_data_out_r[12] , \spi_data_out_r_39__N_1168[12] , \spi_data_out_r_39__N_4835[12] , 
            \spi_data_out_r_39__N_5513[12] , \spi_data_out_r_39__N_4496[12] , 
            \spi_data_out_r_39__N_3818[12] , \spi_data_out_r_39__N_2104[12] , 
            \spi_data_out_r_39__N_1870[12] , \spi_data_out_r_39__N_1402[12] , 
            \spi_data_out_r_39__N_2338[12] , \spi_data_out_r_39__N_5174[12] , 
            \spi_data_out_r_39__N_1636[12] , \spi_data_out_r_39__N_934[12] , 
            \spi_data_out_r_39__N_4157[12] , \spi_data_out_r[13] , \spi_data_out_r_39__N_1168[13] , 
            \spi_data_out_r_39__N_4835[13] , \spi_data_out_r_39__N_5513[13] , 
            \spi_data_out_r_39__N_4496[13] , \spi_data_out_r_39__N_3818[13] , 
            \spi_data_out_r_39__N_2104[13] , \spi_data_out_r_39__N_1870[13] , 
            \spi_data_out_r_39__N_1402[13] , \spi_data_out_r_39__N_2338[13] , 
            \spi_data_out_r_39__N_5174[13] , \spi_data_out_r_39__N_1636[13] , 
            \spi_data_out_r_39__N_934[13] , \spi_data_out_r_39__N_4157[13] , 
            \spi_data_out_r[14] , \spi_data_out_r_39__N_1168[14] , \spi_data_out_r_39__N_4835[14] , 
            \spi_data_out_r_39__N_5513[14] , \spi_data_out_r_39__N_4496[14] , 
            \spi_data_out_r_39__N_3818[14] , \spi_data_out_r_39__N_2104[14] , 
            \spi_data_out_r_39__N_1870[14] , \spi_data_out_r_39__N_1402[14] , 
            \spi_data_out_r_39__N_2338[14] , \spi_data_out_r_39__N_5174[14] , 
            \spi_data_out_r_39__N_1636[14] , \spi_data_out_r_39__N_934[14] , 
            \spi_data_out_r_39__N_4157[14] , \spi_data_out_r[15] , \spi_data_out_r_39__N_1168[15] , 
            \spi_data_out_r_39__N_4835[15] , \spi_data_out_r_39__N_1636[16] , 
            \spi_data_out_r_39__N_5513[15] , \spi_data_out_r_39__N_4496[15] , 
            \spi_data_out_r_39__N_3818[15] , \spi_data_out_r_39__N_2104[15] , 
            \spi_data_out_r_39__N_1870[15] , \spi_data_out_r_39__N_1402[15] , 
            \spi_data_out_r_39__N_2338[15] , \spi_data_out_r_39__N_5174[15] , 
            \spi_data_out_r_39__N_934[16] , \spi_data_out_r_39__N_4157[16] , 
            \spi_data_out_r[17] , \spi_data_out_r_39__N_1168[17] , \spi_data_out_r_39__N_4835[17] , 
            \spi_data_out_r_39__N_5513[17] , \spi_data_out_r_39__N_4496[17] , 
            \spi_data_out_r_39__N_3818[17] , \spi_data_out_r_39__N_2104[17] , 
            \spi_data_out_r_39__N_1870[17] , \spi_data_out_r_39__N_1402[17] , 
            \spi_data_out_r_39__N_2338[17] , \spi_data_out_r_39__N_5174[17] , 
            \spi_data_out_r_39__N_1636[17] , \spi_data_out_r_39__N_934[17] , 
            \spi_data_out_r_39__N_4157[17] , \spi_data_out_r[18] , \spi_data_out_r_39__N_1168[18] , 
            \spi_data_out_r_39__N_4835[18] , \spi_data_out_r_39__N_5513[18] , 
            \spi_data_out_r_39__N_4496[18] , \spi_data_out_r_39__N_3818[18] , 
            \spi_data_out_r_39__N_2104[18] , \spi_data_out_r_39__N_1870[18] , 
            \spi_data_out_r_39__N_1402[18] , \spi_data_out_r_39__N_2338[18] , 
            \spi_data_out_r_39__N_5174[18] , \spi_data_out_r_39__N_1636[18] , 
            \spi_data_out_r_39__N_934[18] , \spi_data_out_r_39__N_4157[18] , 
            \spi_data_out_r[19] , \spi_data_out_r_39__N_1168[19] , \spi_data_out_r_39__N_4835[19] , 
            \spi_data_out_r_39__N_5513[19] , \spi_data_out_r_39__N_4496[19] , 
            \spi_data_out_r_39__N_3818[19] , \spi_data_out_r_39__N_2104[19] , 
            \spi_data_out_r_39__N_1870[19] , \spi_data_out_r_39__N_1402[19] , 
            \spi_data_out_r_39__N_2338[19] , \spi_data_out_r_39__N_5174[19] , 
            \spi_data_out_r_39__N_1636[19] , \spi_data_out_r_39__N_934[19] , 
            \spi_data_out_r_39__N_4157[19] , \spi_data_out_r[20] , \spi_data_out_r_39__N_1168[20] , 
            reset_r, clk_enable_521, n29083, \spi_data_out_r_39__N_4835[20] , 
            \spi_data_out_r_39__N_5513[20] , \spi_data_out_r_39__N_4496[20] , 
            \spi_data_out_r_39__N_3818[20] , \spi_data_out_r_39__N_2104[20] , 
            \spi_data_out_r_39__N_1870[20] , \spi_data_out_r_39__N_1402[20] , 
            \spi_data_out_r_39__N_2338[20] , \spi_data_out_r_39__N_5174[20] , 
            \spi_data_out_r_39__N_1636[20] , \spi_data_out_r_39__N_934[20] , 
            \spi_data_out_r_39__N_4157[20] , \spi_data_out_r[21] , \spi_data_out_r_39__N_1168[21] , 
            \spi_data_out_r_39__N_3818[21] , \spi_data_out_r_39__N_2104[21] , 
            \spi_data_out_r_39__N_1870[21] , \spi_data_out_r_39__N_1402[21] , 
            \spi_data_out_r_39__N_2338[21] , \spi_data_out_r_39__N_5174[21] ) /* synthesis syn_module_defined=1 */ ;
    output \spi_data_out_r[26] ;
    input \spi_data_out_r_39__N_1168[26] ;
    input spi_data_out_r_39__N_1208;
    output [2:0]mode_adj_181;
    input clk;
    input clk_enable_288;
    input n29239;
    input n29762;
    input \spi_data_out_r_39__N_1636[15] ;
    input spi_data_out_r_39__N_1676;
    input \spi_data_out_r_39__N_4835[26] ;
    input spi_data_out_r_39__N_4875;
    input \spi_data_out_r_39__N_5513[26] ;
    input spi_data_out_r_39__N_5553;
    input \spi_data_out_r_39__N_4496[26] ;
    input spi_data_out_r_39__N_4536;
    input \spi_data_out_r_39__N_3818[26] ;
    input spi_data_out_r_39__N_3858;
    input \spi_data_out_r_39__N_2104[26] ;
    input \spi_data_out_r_39__N_1870[26] ;
    input spi_data_out_r_39__N_2144;
    input spi_data_out_r_39__N_1910;
    input \spi_data_out_r_39__N_1402[26] ;
    input spi_data_out_r_39__N_1442;
    input \spi_data_out_r_39__N_2338[26] ;
    input \spi_data_out_r_39__N_5174[26] ;
    input spi_data_out_r_39__N_2378;
    input spi_data_out_r_39__N_5214;
    input \spi_data_out_r_39__N_1636[26] ;
    input \spi_data_out_r_39__N_934[26] ;
    input spi_data_out_r_39__N_974;
    output spi_data_out_r_39__N_5892;
    input \spi_data_out_r_39__N_4157[26] ;
    input spi_data_out_r_39__N_4197;
    input pin_io_out_68;
    output \quad_a[6] ;
    output n28811;
    output \spi_data_out_r[27] ;
    input pin_io_out_69;
    output \quad_b[6] ;
    input \spi_data_out_r_39__N_1168[27] ;
    input \spi_data_out_r_39__N_4835[27] ;
    input \spi_data_out_r_39__N_5513[27] ;
    input \spi_data_out_r_39__N_4835[21] ;
    input \spi_data_out_r_39__N_4496[27] ;
    input \spi_data_out_r_39__N_3818[27] ;
    input \spi_data_out_r_39__N_2104[27] ;
    input \spi_data_out_r_39__N_1870[27] ;
    input \spi_data_out_r_39__N_1402[27] ;
    input \spi_data_out_r_39__N_2338[27] ;
    input \spi_data_out_r_39__N_5174[27] ;
    input \spi_data_out_r_39__N_1636[27] ;
    input \spi_data_out_r_39__N_934[27] ;
    input \spi_data_out_r_39__N_4157[27] ;
    output \spi_data_out_r[28] ;
    input \spi_data_out_r_39__N_1168[28] ;
    output \SLO_buf[0] ;
    output \spi_data_out_r_39__N_5852[0] ;
    input \spi_data_out_r_39__N_6114[0] ;
    input \spi_data_out_r_39__N_4835[28] ;
    input clk_1MHz;
    input clk_1MHz_enable_367;
    input \spi_data_out_r_39__N_5513[28] ;
    input \spi_data_out_r_39__N_934[15] ;
    input \spi_data_out_r_39__N_4157[15] ;
    input \spi_data_out_r_39__N_4496[28] ;
    input \spi_data_out_r_39__N_3818[28] ;
    input \spi_data_out_r_39__N_2104[28] ;
    input \spi_data_out_r_39__N_1870[28] ;
    input \spi_data_out_r_39__N_1402[28] ;
    input \spi_data_out_r_39__N_2338[28] ;
    input \spi_data_out_r_39__N_5174[28] ;
    input \spi_data_out_r_39__N_1636[21] ;
    input \spi_data_out_r_39__N_934[21] ;
    input \spi_data_out_r_39__N_4157[21] ;
    input \spi_data_out_r_39__N_1636[28] ;
    output \spi_data_out_r[22] ;
    input \spi_data_out_r_39__N_1168[22] ;
    input \spi_data_out_r_39__N_4835[22] ;
    input \spi_data_out_r_39__N_5513[22] ;
    input \spi_data_out_r_39__N_934[28] ;
    input \spi_data_out_r_39__N_4157[28] ;
    output \spi_data_out_r[29] ;
    input \spi_data_out_r_39__N_4496[22] ;
    input \spi_data_out_r_39__N_1168[29] ;
    input \spi_data_out_r_39__N_4835[29] ;
    input \spi_data_out_r_39__N_5513[29] ;
    input \spi_data_out_r_39__N_4496[29] ;
    input \spi_data_out_r_39__N_3818[29] ;
    input \spi_data_out_r_39__N_3818[22] ;
    input \spi_data_out_r_39__N_2104[29] ;
    input \spi_data_out_r_39__N_1870[29] ;
    input \spi_data_out_r_39__N_2104[22] ;
    input \spi_data_out_r_39__N_1870[22] ;
    input \spi_data_out_r_39__N_1402[22] ;
    input \spi_data_out_r_39__N_1402[29] ;
    input \spi_data_out_r_39__N_2338[29] ;
    input \spi_data_out_r_39__N_5174[29] ;
    input \spi_data_out_r_39__N_1636[29] ;
    input \spi_data_out_r_39__N_2338[22] ;
    input \spi_data_out_r_39__N_5174[22] ;
    input \spi_data_out_r_39__N_934[29] ;
    input n29087;
    input \spi_data_out_r_39__N_4157[29] ;
    input \spi_data_out_r_39__N_1636[22] ;
    output \spi_data_out_r[30] ;
    input \spi_data_out_r_39__N_1168[30] ;
    input \spi_data_out_r_39__N_934[22] ;
    input \spi_data_out_r_39__N_4835[30] ;
    input \spi_data_out_r_39__N_5513[30] ;
    input \spi_data_out_r_39__N_4157[22] ;
    input \spi_data_out_r_39__N_4496[30] ;
    output \spi_data_out_r[23] ;
    input \spi_data_out_r_39__N_3818[30] ;
    output digital_output_r;
    input clk_enable_198;
    input \spi_data_r[0] ;
    input \spi_data_out_r_39__N_1168[23] ;
    input \spi_data_out_r_39__N_2104[30] ;
    input \spi_data_out_r_39__N_1870[30] ;
    input \spi_data_out_r_39__N_1402[30] ;
    input \spi_data_out_r_39__N_2338[30] ;
    input \spi_data_out_r_39__N_5174[30] ;
    input \spi_data_out_r_39__N_1636[30] ;
    input \spi_data_out_r_39__N_934[30] ;
    input \spi_data_out_r_39__N_4157[30] ;
    output \spi_data_out_r[31] ;
    input \spi_data_out_r_39__N_4835[23] ;
    input \spi_data_out_r_39__N_1168[31] ;
    input \spi_data_out_r_39__N_5513[23] ;
    output \spi_data_out_r[16] ;
    input \spi_data_out_r_39__N_1168[16] ;
    input \spi_data_out_r_39__N_4496[23] ;
    input \spi_data_out_r_39__N_4835[31] ;
    input \spi_data_out_r_39__N_3818[23] ;
    input \spi_data_out_r_39__N_5513[31] ;
    input \spi_data_out_r_39__N_4496[31] ;
    output n19401;
    input resetn_c;
    input \spi_data_out_r_39__N_3818[31] ;
    input \spi_data_out_r_39__N_2104[31] ;
    input \spi_data_out_r_39__N_1870[31] ;
    input \spi_data_out_r_39__N_1402[31] ;
    input \spi_data_out_r_39__N_2338[31] ;
    input \spi_data_out_r_39__N_5174[31] ;
    input \spi_data_out_r_39__N_1636[31] ;
    input \spi_data_out_r_39__N_934[31] ;
    input \spi_data_out_r_39__N_4157[31] ;
    input \spi_data_out_r_39__N_4835[32] ;
    output \spi_data_out_r[32] ;
    input \spi_data_out_r_39__N_3818[32] ;
    input \spi_data_out_r_39__N_5174[32] ;
    input \spi_data_out_r_39__N_4496[32] ;
    input \spi_data_out_r_39__N_4157[32] ;
    input \spi_data_out_r_39__N_5513[32] ;
    input \spi_data_out_r_39__N_4835[33] ;
    output \spi_data_out_r[33] ;
    input \spi_data_out_r_39__N_3818[33] ;
    input \spi_data_out_r_39__N_5174[33] ;
    input \spi_data_out_r_39__N_4496[33] ;
    input \spi_data_out_r_39__N_4157[33] ;
    input \spi_data_out_r_39__N_5513[33] ;
    input \spi_data_out_r_39__N_4835[34] ;
    output \spi_data_out_r[34] ;
    input \spi_data_out_r_39__N_3818[34] ;
    input \spi_data_out_r_39__N_5174[34] ;
    input \spi_data_out_r_39__N_4496[34] ;
    input \spi_data_out_r_39__N_4157[34] ;
    input \spi_data_out_r_39__N_2104[23] ;
    input \spi_data_out_r_39__N_1870[23] ;
    input \spi_data_out_r_39__N_5513[34] ;
    input \spi_data_out_r_39__N_4835[35] ;
    output \spi_data_out_r[35] ;
    input \spi_data_out_r_39__N_3818[35] ;
    input \spi_data_out_r_39__N_5174[35] ;
    input \spi_data_out_r_39__N_4496[35] ;
    input \spi_data_out_r_39__N_4157[35] ;
    input \spi_data_out_r_39__N_5513[35] ;
    input \spi_data_out_r_39__N_4835[36] ;
    output \spi_data_out_r[36] ;
    input \spi_data_out_r_39__N_3818[36] ;
    input \spi_data_out_r_39__N_5174[36] ;
    input \spi_data_out_r_39__N_4496[36] ;
    input \spi_data_out_r_39__N_4157[36] ;
    input \spi_data_out_r_39__N_5513[36] ;
    input \spi_data_out_r_39__N_4835[37] ;
    output \spi_data_out_r[37] ;
    input \spi_data_out_r_39__N_1402[23] ;
    input \spi_data_out_r_39__N_3818[37] ;
    input \spi_data_out_r_39__N_5174[37] ;
    input \spi_data_out_r_39__N_4496[37] ;
    input \spi_data_out_r_39__N_4157[37] ;
    input \spi_data_out_r_39__N_2338[23] ;
    input \spi_data_out_r_39__N_5174[23] ;
    input \spi_data_out_r_39__N_5513[37] ;
    input \spi_data_out_r_39__N_4835[38] ;
    output \spi_data_out_r[38] ;
    input \spi_data_out_r_39__N_3818[38] ;
    input \spi_data_out_r_39__N_1636[23] ;
    input \spi_data_out_r_39__N_5174[38] ;
    input \spi_data_out_r_39__N_4496[38] ;
    input \spi_data_out_r_39__N_4157[38] ;
    input \spi_data_out_r_39__N_934[23] ;
    input \spi_data_out_r_39__N_4157[23] ;
    input \spi_data_out_r_39__N_5513[38] ;
    input \spi_data_out_r_39__N_4835[39] ;
    output \spi_data_out_r[39] ;
    input \spi_data_out_r_39__N_3818[39] ;
    input \spi_data_out_r_39__N_5174[39] ;
    input \spi_data_out_r_39__N_4496[39] ;
    input \spi_data_out_r_39__N_4157[39] ;
    input \spi_data_out_r_39__N_5513[39] ;
    output \spi_data_out_r[24] ;
    input \spi_data_out_r_39__N_1168[24] ;
    input \spi_data_out_r_39__N_4835[24] ;
    input \spi_data_out_r_39__N_5513[24] ;
    input \spi_data_out_r_39__N_4496[24] ;
    input n29267;
    input mode;
    input n29191;
    output n29153;
    input \spi_data_out_r_39__N_3818[24] ;
    output n29195;
    input \spi_data_out_r_39__N_2104[24] ;
    input \spi_data_out_r_39__N_1870[24] ;
    input n29293;
    input \cs_decoded[12] ;
    output n8652;
    output n1;
    output n8651;
    output n1_adj_171;
    input \spi_data_out_r_39__N_5513[21] ;
    input \spi_data_out_r_39__N_1402[24] ;
    input \spi_data_out_r_39__N_2338[24] ;
    input \spi_data_out_r_39__N_5174[24] ;
    input \spi_data_out_r_39__N_1636[24] ;
    input \spi_data_out_r_39__N_934[24] ;
    input \spi_data_out_r_39__N_4157[24] ;
    output \spi_data_out_r[25] ;
    input \spi_data_out_r_39__N_1168[25] ;
    input \spi_data_out_r_39__N_4835[25] ;
    input \spi_data_out_r_39__N_5513[25] ;
    input \spi_data_out_r_39__N_4496[25] ;
    input \spi_data_out_r_39__N_3818[25] ;
    input \spi_data_out_r_39__N_2104[25] ;
    input \spi_data_out_r_39__N_1870[25] ;
    input \spi_data_out_r_39__N_1402[25] ;
    input \spi_data_out_r_39__N_2338[25] ;
    input \spi_data_out_r_39__N_5174[25] ;
    input GND_net;
    input \spi_data_out_r_39__N_1636[25] ;
    input \spi_data_out_r_39__N_934[25] ;
    input \spi_data_out_r_39__N_4157[25] ;
    input \spi_data_r[2] ;
    input \spi_data_r[1] ;
    input \spi_data_out_r_39__N_4835[16] ;
    input \spi_data_out_r_39__N_2856[2] ;
    input clear_intrpt;
    output n13;
    input \spi_data_out_r_39__N_1402[2] ;
    output n4;
    output \SLO_buf[1] ;
    output \SLO_buf[2] ;
    output \SLO_buf[3] ;
    output \SLO_buf[4] ;
    output \SLO_buf[5] ;
    output \SLO_buf[6] ;
    output \SLO_buf[7] ;
    output \SLO_buf[8] ;
    output \SLO_buf[9] ;
    output \SLO_buf[10] ;
    output \SLO_buf[11] ;
    output \SLO_buf[12] ;
    output \SLO_buf[13] ;
    output \SLO_buf[14] ;
    output \SLO_buf[15] ;
    output \SLO_buf[16] ;
    output \SLO_buf[17] ;
    output \SLO_buf[18] ;
    output \SLO_buf[19] ;
    output \SLO_buf[20] ;
    output \SLO_buf[21] ;
    output \SLO_buf[22] ;
    output \SLO_buf[23] ;
    output \SLO_buf[24] ;
    output \SLO_buf[25] ;
    output \SLO_buf[26] ;
    output \SLO_buf[27] ;
    output \SLO_buf[28] ;
    output \SLO_buf[29] ;
    input \spi_data_out_r_39__N_5513[16] ;
    input \spi_data_out_r_39__N_6114[1] ;
    output \spi_data_out_r_39__N_5852[2] ;
    input \spi_data_out_r_39__N_6114[2] ;
    input \spi_data_out_r_39__N_6114[3] ;
    input \spi_data_out_r_39__N_6114[4] ;
    input \spi_data_out_r_39__N_6114[5] ;
    input \spi_data_out_r_39__N_6114[6] ;
    input \spi_data_out_r_39__N_6114[7] ;
    input \spi_data_out_r_39__N_6114[8] ;
    input \spi_data_out_r_39__N_6114[9] ;
    input \spi_data_out_r_39__N_6114[10] ;
    input \spi_data_out_r_39__N_6114[11] ;
    input \spi_data_out_r_39__N_6114[12] ;
    input \spi_data_out_r_39__N_6114[13] ;
    input \spi_data_out_r_39__N_6114[14] ;
    input \spi_data_out_r_39__N_6114[15] ;
    input n29076;
    input \spi_data_out_r_39__N_6114[32] ;
    input \spi_data_out_r_39__N_6114[33] ;
    input \spi_data_out_r_39__N_6114[34] ;
    input \spi_data_out_r_39__N_6114[35] ;
    input \spi_data_out_r_39__N_4496[16] ;
    input \spi_data_out_r_39__N_2338[2] ;
    output n8;
    input \spi_data_out_r_39__N_2998[2] ;
    input clear_intrpt_adj_172;
    output n15;
    input \spi_data_out_r_39__N_2714[2] ;
    input clear_intrpt_adj_173;
    output n11;
    input \spi_data_out_r_39__N_4835[2] ;
    output n19;
    input \spi_data_out_r_39__N_3818[16] ;
    input \spi_data_out_r_39__N_4157[0] ;
    output n17;
    input \spi_data_out_r_39__N_1168[0] ;
    output n3;
    input \spi_data_out_r_39__N_5174[0] ;
    output n20;
    input \spi_data_out_r_39__N_2998[0] ;
    output n15_adj_174;
    input \spi_data_out_r_39__N_934[0] ;
    output n2;
    input \spi_data_out_r_39__N_5513[0] ;
    output n21;
    input \spi_data_out_r_39__N_1402[0] ;
    output n4_adj_175;
    input \spi_data_out_r_39__N_2714[0] ;
    output n11_adj_176;
    output \spi_data_out_r[1] ;
    input \spi_data_out_r_39__N_2643[1] ;
    input \spi_data_out_r_39__N_2856[1] ;
    input clear_intrpt_adj_177;
    input \spi_data_out_r_39__N_934[1] ;
    input \spi_data_out_r_39__N_4157[1] ;
    input \spi_data_out_r_39__N_1168[1] ;
    input \spi_data_out_r_39__N_2927[1] ;
    input \spi_data_out_r_39__N_2785[1] ;
    input clear_intrpt_adj_178;
    input clear_intrpt_adj_179;
    input \spi_data_out_r_39__N_1402[1] ;
    input \spi_data_out_r_39__N_5174[1] ;
    input \spi_data_out_r_39__N_3818[1] ;
    input \spi_data_out_r_39__N_2338[1] ;
    input \spi_data_out_r_39__N_4496[21] ;
    input \spi_data_out_r_39__N_4496[1] ;
    input \spi_data_out_r_39__N_1870[1] ;
    input \spi_data_out_r_39__N_2998[1] ;
    input \spi_data_out_r_39__N_2104[1] ;
    input \spi_data_out_r_39__N_2572[1] ;
    input clear_intrpt_adj_180;
    input \spi_data_out_r_39__N_4835[1] ;
    input \spi_data_out_r_39__N_5513[1] ;
    input \spi_data_out_r_39__N_1636[1] ;
    input \spi_data_out_r_39__N_2714[1] ;
    output \spi_data_out_r[3] ;
    input \spi_data_out_r_39__N_1168[3] ;
    input \spi_data_out_r_39__N_4835[3] ;
    input \spi_data_out_r_39__N_5513[3] ;
    input \spi_data_out_r_39__N_4496[3] ;
    input \spi_data_out_r_39__N_3818[3] ;
    input \spi_data_out_r_39__N_2104[3] ;
    input \spi_data_out_r_39__N_1870[3] ;
    input \spi_data_out_r_39__N_1402[3] ;
    input \spi_data_out_r_39__N_2338[3] ;
    input \spi_data_out_r_39__N_5174[3] ;
    input \spi_data_out_r_39__N_1636[3] ;
    input \spi_data_out_r_39__N_934[3] ;
    input \spi_data_out_r_39__N_4157[3] ;
    output \spi_data_out_r[4] ;
    input \spi_data_out_r_39__N_1168[4] ;
    input \spi_data_out_r_39__N_4835[4] ;
    input \spi_data_out_r_39__N_5513[4] ;
    input \spi_data_out_r_39__N_4496[4] ;
    input \spi_data_out_r_39__N_2104[16] ;
    input \spi_data_out_r_39__N_1870[16] ;
    input \spi_data_out_r_39__N_3818[4] ;
    input \spi_data_out_r_39__N_2104[4] ;
    input \spi_data_out_r_39__N_1870[4] ;
    input \spi_data_out_r_39__N_1402[16] ;
    input \spi_data_out_r_39__N_1402[4] ;
    input \spi_data_out_r_39__N_2338[4] ;
    input \spi_data_out_r_39__N_5174[4] ;
    input \spi_data_out_r_39__N_1636[4] ;
    input \spi_data_out_r_39__N_934[4] ;
    input \spi_data_out_r_39__N_4157[4] ;
    output \spi_data_out_r[5] ;
    input \spi_data_out_r_39__N_1168[5] ;
    input \spi_data_out_r_39__N_4835[5] ;
    input \spi_data_out_r_39__N_5513[5] ;
    input \spi_data_out_r_39__N_4496[5] ;
    input \spi_data_out_r_39__N_3818[5] ;
    input \spi_data_out_r_39__N_2104[5] ;
    input \spi_data_out_r_39__N_1870[5] ;
    input \spi_data_out_r_39__N_1402[5] ;
    input \spi_data_out_r_39__N_2338[5] ;
    input \spi_data_out_r_39__N_5174[5] ;
    input \spi_data_out_r_39__N_1636[5] ;
    input \spi_data_out_r_39__N_934[5] ;
    input \spi_data_out_r_39__N_4157[5] ;
    output \spi_data_out_r[6] ;
    input \spi_data_out_r_39__N_1168[6] ;
    input \spi_data_out_r_39__N_4835[6] ;
    input \spi_data_out_r_39__N_5513[6] ;
    input \spi_data_out_r_39__N_4496[6] ;
    input \spi_data_out_r_39__N_3818[6] ;
    input \spi_data_out_r_39__N_2104[6] ;
    input \spi_data_out_r_39__N_1870[6] ;
    input \spi_data_out_r_39__N_1402[6] ;
    input \spi_data_out_r_39__N_2338[6] ;
    input \spi_data_out_r_39__N_5174[6] ;
    input \spi_data_out_r_39__N_1636[6] ;
    input \spi_data_out_r_39__N_934[6] ;
    input \spi_data_out_r_39__N_4157[6] ;
    output \spi_data_out_r[7] ;
    input \spi_data_out_r_39__N_1168[7] ;
    input \spi_data_out_r_39__N_4835[7] ;
    input \spi_data_out_r_39__N_5513[7] ;
    input \spi_data_out_r_39__N_4496[7] ;
    input \spi_data_out_r_39__N_3818[7] ;
    input \spi_data_out_r_39__N_2104[7] ;
    input \spi_data_out_r_39__N_1870[7] ;
    input \spi_data_out_r_39__N_1402[7] ;
    input \spi_data_out_r_39__N_2338[7] ;
    input \spi_data_out_r_39__N_5174[7] ;
    input \spi_data_out_r_39__N_1636[7] ;
    input \spi_data_out_r_39__N_934[7] ;
    input \spi_data_out_r_39__N_4157[7] ;
    output \spi_data_out_r[8] ;
    input \spi_data_out_r_39__N_1168[8] ;
    input \spi_data_out_r_39__N_4835[8] ;
    input \spi_data_out_r_39__N_5513[8] ;
    input \spi_data_out_r_39__N_4496[8] ;
    input \spi_data_out_r_39__N_3818[8] ;
    input \spi_data_out_r_39__N_2104[8] ;
    input \spi_data_out_r_39__N_1870[8] ;
    input \spi_data_out_r_39__N_1402[8] ;
    input \spi_data_out_r_39__N_2338[8] ;
    input \spi_data_out_r_39__N_5174[8] ;
    input \spi_data_out_r_39__N_1636[8] ;
    input \spi_data_out_r_39__N_934[8] ;
    input \spi_data_out_r_39__N_4157[8] ;
    output \spi_data_out_r[9] ;
    input \spi_data_out_r_39__N_1168[9] ;
    input \spi_data_out_r_39__N_4835[9] ;
    input \spi_data_out_r_39__N_5513[9] ;
    input \spi_data_out_r_39__N_4496[9] ;
    input \spi_data_out_r_39__N_3818[9] ;
    input \spi_data_out_r_39__N_2104[9] ;
    input \spi_data_out_r_39__N_1870[9] ;
    input \spi_data_out_r_39__N_1402[9] ;
    input \spi_data_out_r_39__N_2338[9] ;
    input \spi_data_out_r_39__N_5174[9] ;
    input \spi_data_out_r_39__N_1636[9] ;
    input \spi_data_out_r_39__N_2338[16] ;
    input \spi_data_out_r_39__N_5174[16] ;
    input \spi_data_out_r_39__N_934[9] ;
    input \spi_data_out_r_39__N_4157[9] ;
    output \spi_data_out_r[10] ;
    input \spi_data_out_r_39__N_1168[10] ;
    input \spi_data_out_r_39__N_4835[10] ;
    input \spi_data_out_r_39__N_5513[10] ;
    input \spi_data_out_r_39__N_4496[10] ;
    input \spi_data_out_r_39__N_3818[10] ;
    input \spi_data_out_r_39__N_2104[10] ;
    input \spi_data_out_r_39__N_1870[10] ;
    input \spi_data_out_r_39__N_1402[10] ;
    input \spi_data_out_r_39__N_2338[10] ;
    input \spi_data_out_r_39__N_5174[10] ;
    input \spi_data_out_r_39__N_1636[10] ;
    input \spi_data_out_r_39__N_934[10] ;
    input \spi_data_out_r_39__N_4157[10] ;
    output \spi_data_out_r[11] ;
    input \spi_data_out_r_39__N_1168[11] ;
    input \spi_data_out_r_39__N_4835[11] ;
    input \spi_data_out_r_39__N_5513[11] ;
    input \spi_data_out_r_39__N_4496[11] ;
    input \spi_data_out_r_39__N_3818[11] ;
    input \spi_data_out_r_39__N_2104[11] ;
    input \spi_data_out_r_39__N_1870[11] ;
    input \spi_data_out_r_39__N_1402[11] ;
    input \spi_data_out_r_39__N_2338[11] ;
    input \spi_data_out_r_39__N_5174[11] ;
    input \spi_data_out_r_39__N_1636[11] ;
    input \spi_data_out_r_39__N_934[11] ;
    input \spi_data_out_r_39__N_4157[11] ;
    output \spi_data_out_r[12] ;
    input \spi_data_out_r_39__N_1168[12] ;
    input \spi_data_out_r_39__N_4835[12] ;
    input \spi_data_out_r_39__N_5513[12] ;
    input \spi_data_out_r_39__N_4496[12] ;
    input \spi_data_out_r_39__N_3818[12] ;
    input \spi_data_out_r_39__N_2104[12] ;
    input \spi_data_out_r_39__N_1870[12] ;
    input \spi_data_out_r_39__N_1402[12] ;
    input \spi_data_out_r_39__N_2338[12] ;
    input \spi_data_out_r_39__N_5174[12] ;
    input \spi_data_out_r_39__N_1636[12] ;
    input \spi_data_out_r_39__N_934[12] ;
    input \spi_data_out_r_39__N_4157[12] ;
    output \spi_data_out_r[13] ;
    input \spi_data_out_r_39__N_1168[13] ;
    input \spi_data_out_r_39__N_4835[13] ;
    input \spi_data_out_r_39__N_5513[13] ;
    input \spi_data_out_r_39__N_4496[13] ;
    input \spi_data_out_r_39__N_3818[13] ;
    input \spi_data_out_r_39__N_2104[13] ;
    input \spi_data_out_r_39__N_1870[13] ;
    input \spi_data_out_r_39__N_1402[13] ;
    input \spi_data_out_r_39__N_2338[13] ;
    input \spi_data_out_r_39__N_5174[13] ;
    input \spi_data_out_r_39__N_1636[13] ;
    input \spi_data_out_r_39__N_934[13] ;
    input \spi_data_out_r_39__N_4157[13] ;
    output \spi_data_out_r[14] ;
    input \spi_data_out_r_39__N_1168[14] ;
    input \spi_data_out_r_39__N_4835[14] ;
    input \spi_data_out_r_39__N_5513[14] ;
    input \spi_data_out_r_39__N_4496[14] ;
    input \spi_data_out_r_39__N_3818[14] ;
    input \spi_data_out_r_39__N_2104[14] ;
    input \spi_data_out_r_39__N_1870[14] ;
    input \spi_data_out_r_39__N_1402[14] ;
    input \spi_data_out_r_39__N_2338[14] ;
    input \spi_data_out_r_39__N_5174[14] ;
    input \spi_data_out_r_39__N_1636[14] ;
    input \spi_data_out_r_39__N_934[14] ;
    input \spi_data_out_r_39__N_4157[14] ;
    output \spi_data_out_r[15] ;
    input \spi_data_out_r_39__N_1168[15] ;
    input \spi_data_out_r_39__N_4835[15] ;
    input \spi_data_out_r_39__N_1636[16] ;
    input \spi_data_out_r_39__N_5513[15] ;
    input \spi_data_out_r_39__N_4496[15] ;
    input \spi_data_out_r_39__N_3818[15] ;
    input \spi_data_out_r_39__N_2104[15] ;
    input \spi_data_out_r_39__N_1870[15] ;
    input \spi_data_out_r_39__N_1402[15] ;
    input \spi_data_out_r_39__N_2338[15] ;
    input \spi_data_out_r_39__N_5174[15] ;
    input \spi_data_out_r_39__N_934[16] ;
    input \spi_data_out_r_39__N_4157[16] ;
    output \spi_data_out_r[17] ;
    input \spi_data_out_r_39__N_1168[17] ;
    input \spi_data_out_r_39__N_4835[17] ;
    input \spi_data_out_r_39__N_5513[17] ;
    input \spi_data_out_r_39__N_4496[17] ;
    input \spi_data_out_r_39__N_3818[17] ;
    input \spi_data_out_r_39__N_2104[17] ;
    input \spi_data_out_r_39__N_1870[17] ;
    input \spi_data_out_r_39__N_1402[17] ;
    input \spi_data_out_r_39__N_2338[17] ;
    input \spi_data_out_r_39__N_5174[17] ;
    input \spi_data_out_r_39__N_1636[17] ;
    input \spi_data_out_r_39__N_934[17] ;
    input \spi_data_out_r_39__N_4157[17] ;
    output \spi_data_out_r[18] ;
    input \spi_data_out_r_39__N_1168[18] ;
    input \spi_data_out_r_39__N_4835[18] ;
    input \spi_data_out_r_39__N_5513[18] ;
    input \spi_data_out_r_39__N_4496[18] ;
    input \spi_data_out_r_39__N_3818[18] ;
    input \spi_data_out_r_39__N_2104[18] ;
    input \spi_data_out_r_39__N_1870[18] ;
    input \spi_data_out_r_39__N_1402[18] ;
    input \spi_data_out_r_39__N_2338[18] ;
    input \spi_data_out_r_39__N_5174[18] ;
    input \spi_data_out_r_39__N_1636[18] ;
    input \spi_data_out_r_39__N_934[18] ;
    input \spi_data_out_r_39__N_4157[18] ;
    output \spi_data_out_r[19] ;
    input \spi_data_out_r_39__N_1168[19] ;
    input \spi_data_out_r_39__N_4835[19] ;
    input \spi_data_out_r_39__N_5513[19] ;
    input \spi_data_out_r_39__N_4496[19] ;
    input \spi_data_out_r_39__N_3818[19] ;
    input \spi_data_out_r_39__N_2104[19] ;
    input \spi_data_out_r_39__N_1870[19] ;
    input \spi_data_out_r_39__N_1402[19] ;
    input \spi_data_out_r_39__N_2338[19] ;
    input \spi_data_out_r_39__N_5174[19] ;
    input \spi_data_out_r_39__N_1636[19] ;
    input \spi_data_out_r_39__N_934[19] ;
    input \spi_data_out_r_39__N_4157[19] ;
    output \spi_data_out_r[20] ;
    input \spi_data_out_r_39__N_1168[20] ;
    output reset_r;
    input clk_enable_521;
    input n29083;
    input \spi_data_out_r_39__N_4835[20] ;
    input \spi_data_out_r_39__N_5513[20] ;
    input \spi_data_out_r_39__N_4496[20] ;
    input \spi_data_out_r_39__N_3818[20] ;
    input \spi_data_out_r_39__N_2104[20] ;
    input \spi_data_out_r_39__N_1870[20] ;
    input \spi_data_out_r_39__N_1402[20] ;
    input \spi_data_out_r_39__N_2338[20] ;
    input \spi_data_out_r_39__N_5174[20] ;
    input \spi_data_out_r_39__N_1636[20] ;
    input \spi_data_out_r_39__N_934[20] ;
    input \spi_data_out_r_39__N_4157[20] ;
    output \spi_data_out_r[21] ;
    input \spi_data_out_r_39__N_1168[21] ;
    input \spi_data_out_r_39__N_3818[21] ;
    input \spi_data_out_r_39__N_2104[21] ;
    input \spi_data_out_r_39__N_1870[21] ;
    input \spi_data_out_r_39__N_1402[21] ;
    input \spi_data_out_r_39__N_2338[21] ;
    input \spi_data_out_r_39__N_5174[21] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire MA_Temp_N_5969 /* synthesis is_inv_clock=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    wire clk_1MHz_derived_322 /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz_derived_322 */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire MA_Temp /* synthesis is_clock=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(57[5:12])
    
    wire n3_c, n26, n22, n21_c, n18, n24, n18_adj_6759, n4_c, 
        n5, n16, n17_c, n20_c, n5_adj_6760;
    wire [39:0]spi_data_out_r_39__N_5852;
    
    wire n3_adj_6761, n26_adj_6762, n22_adj_6763, n21_adj_6764, n18_adj_6765, 
        n24_adj_6766, n18_adj_6767, n4_adj_6768, n16_adj_6769, n17_adj_6770, 
        n16_adj_6771, n17_adj_6772, n22_adj_6773, n20_adj_6774, n5_adj_6775, 
        n3_adj_6776, n26_adj_6777, n22_adj_6778, n21_adj_6779, n18_adj_6780, 
        n24_adj_6781, n18_adj_6782, n4_adj_6783;
    wire [51:0]SLO;   // c:/s_links/sources/slot_cards/stepper.v(63[12:15])
    
    wire clk_1MHz_derived_322_enable_20, n16_adj_6784, n17_adj_6785;
    wire [11:0]Cnt_NSL;   // c:/s_links/sources/slot_cards/stepper.v(61[12:19])
    wire [11:0]n1290;
    wire [7:0]Cnt;   // c:/s_links/sources/slot_cards/stepper.v(62[11:14])
    
    wire clk_1MHz_enable_374;
    wire [7:0]n199;
    
    wire n16_adj_6786, n17_adj_6787, n20_adj_6788, n5_adj_6789, n5_adj_6790, 
        n3_adj_6791, n26_adj_6792, n22_adj_6793, n21_adj_6794, n18_adj_6795, 
        n24_adj_6796, n18_adj_6797, n4_adj_6798, n16_adj_6799, n17_adj_6800, 
        n3_adj_6801, n26_adj_6802, n22_adj_6803, n21_adj_6804, n18_adj_6805, 
        n24_adj_6806, n18_adj_6807, n4_adj_6808, n16_adj_6809, n17_adj_6810, 
        n20_adj_6811, n5_adj_6812, n20_adj_6813, n5_adj_6814, n28796, 
        n28795, n19545, n28797, n3_adj_6815, n26_adj_6816, n22_adj_6817, 
        n21_adj_6818, n18_adj_6819, n24_adj_6820, n18_adj_6821, n4_adj_6822, 
        n16_adj_6823, n17_adj_6824, n3_adj_6825, n26_adj_6826, n22_adj_6827, 
        n21_adj_6828, n20_adj_6829, n5_adj_6830, n18_adj_6831, n24_adj_6832, 
        n18_adj_6833, n4_adj_6834, n3_adj_6835, n26_adj_6836, n22_adj_6837, 
        n21_adj_6838, n16_adj_6839, n17_adj_6840, n3_adj_6841, n26_adj_6842, 
        n22_adj_6843, n21_adj_6844, n18_adj_6845, n24_adj_6846, n18_adj_6847, 
        n4_adj_6848, n16_adj_6849, n17_adj_6850, n20_adj_6851, n5_adj_6852, 
        n20_adj_6853, n5_adj_6854, n19439, clk_1MHz_enable_377, n12, 
        n8_c, n10, n21_adj_6855, n12_adj_6856, n8_adj_6857, n10_adj_6858, 
        n21_adj_6859, n12_adj_6860, n8_adj_6861, n10_adj_6862, n21_adj_6863, 
        n12_adj_6864, n8_adj_6865, n10_adj_6866, n21_adj_6867, n12_adj_6868, 
        n8_adj_6869, n10_adj_6870, n21_adj_6871, n12_adj_6872, n8_adj_6873, 
        n10_adj_6874, n21_adj_6875, n12_adj_6876, n8_adj_6877, n10_adj_6878, 
        n21_adj_6879, n12_adj_6880, n8_adj_6881, n10_adj_6882, n21_adj_6883, 
        n29271, n29192, n11795, n3_adj_6884, n26_adj_6885, n22_adj_6886, 
        n21_adj_6887, n18_adj_6888, n24_adj_6889, n18_adj_6890, n4_adj_6891, 
        n16_adj_6892, n17_adj_6893, n20_adj_6894, n5_adj_6895, n29275, 
        n27387, n29156, n29277, MA_Temp_N_5983, n13378, NSL, clk_1MHz_derived_322_enable_46, 
        n21_adj_6897, n3_adj_6898, n26_adj_6899, n22_adj_6900, n21_adj_6901, 
        n18_adj_6902, n24_adj_6903, n18_adj_6904, n4_adj_6905, n16_adj_6906, 
        n17_adj_6907, n20_adj_6908, n5_adj_6909, n25044, n25043, n25042, 
        n25041, n25040, clk_1MHz_enable_247, NSL_N_6180, n25039, n25038;
    wire [31:0]n153;
    
    wire n18_adj_6910, n24_adj_6911, n18_adj_6912, n4_adj_6913, n16_adj_6914, 
        n17_adj_6915;
    wire [51:0]SLO_buf;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire n4_adj_6918, n25037, n25036, n19465, n20_adj_6921, n5_adj_6922, 
        n25035, n28794, n27, n40, n36, n28, n31, n38, n4_adj_6931, 
        n22_adj_6932, n30, n19_adj_6933, n8_adj_6936, n34, n24_adj_6937, 
        n15_adj_6938, n18_adj_6939, n26_adj_6940, n11_adj_6941, n3_adj_6943, 
        n26_adj_6944, n22_adj_6945, n21_adj_6946, n18_adj_6947, n24_adj_6948, 
        n18_adj_6949, n4_adj_6950, n16_adj_6951, n17_adj_6952, MA_Temp_N_5972, 
        n20_adj_6953, n5_adj_6954, n3_adj_6955, n26_adj_6956, n22_adj_6957, 
        n21_adj_6958, n18_adj_6959, n24_adj_6960, n18_adj_6961, n4_adj_6962, 
        n16_adj_6963, n17_adj_6964, n20_adj_6965, n5_adj_6966, n3_adj_6967, 
        n26_adj_6968, n22_adj_6969, n21_adj_6970, n18_adj_6971, n24_adj_6972, 
        n18_adj_6973, n4_adj_6974, n16_adj_6975, n17_adj_6976, n20_adj_6977, 
        n5_adj_6978, n3_adj_6979, n26_adj_6980, n22_adj_6981, n21_adj_6982, 
        n18_adj_6983, n24_adj_6984, n18_adj_6985, n4_adj_6986, n16_adj_6987, 
        n17_adj_6988, n20_adj_6989, n5_adj_6990, n3_adj_6991, n26_adj_6992, 
        n22_adj_6993, n21_adj_6994, n18_adj_6995, n24_adj_6996, n18_adj_6997, 
        n4_adj_6998, n16_adj_6999, n17_adj_7000, n20_adj_7001, n5_adj_7002, 
        n3_adj_7003, n26_adj_7004, n22_adj_7005, n21_adj_7006, n18_adj_7007, 
        n24_adj_7008, n18_adj_7009, n4_adj_7010, n16_adj_7011, n17_adj_7012, 
        n20_adj_7013, n5_adj_7014, n3_adj_7015, n26_adj_7016, n22_adj_7017, 
        n21_adj_7018, n18_adj_7019, n24_adj_7020, n18_adj_7021, n4_adj_7022, 
        n16_adj_7023, n17_adj_7024, n20_adj_7025, n5_adj_7026, n3_adj_7027, 
        n26_adj_7028, n22_adj_7029, n21_adj_7030, n18_adj_7031, n24_adj_7032, 
        n18_adj_7033, n4_adj_7034, n16_adj_7035, n17_adj_7036, n20_adj_7037, 
        n5_adj_7038, n3_adj_7039, n26_adj_7040, n22_adj_7041, n21_adj_7042, 
        n18_adj_7043, n24_adj_7044, n18_adj_7045, n4_adj_7046, n16_adj_7047, 
        n17_adj_7048, n20_adj_7049, n5_adj_7050, n3_adj_7051, n26_adj_7052, 
        n22_adj_7053, n21_adj_7054, n18_adj_7055, n24_adj_7056, n18_adj_7057, 
        n4_adj_7058, n16_adj_7059, n17_adj_7060, n20_adj_7061, n5_adj_7062, 
        n3_adj_7063, n26_adj_7064, n22_adj_7065, n21_adj_7066, n18_adj_7067, 
        n24_adj_7068, n18_adj_7069, n4_adj_7070, n16_adj_7071, n17_adj_7072, 
        n20_adj_7073, n5_adj_7074, n3_adj_7075, n26_adj_7076, n22_adj_7077, 
        n21_adj_7078, n18_adj_7079, n24_adj_7080, n18_adj_7081, n4_adj_7082, 
        n16_adj_7083, n17_adj_7084, n20_adj_7085, n5_adj_7086, n3_adj_7087, 
        n26_adj_7088, n22_adj_7089, n21_adj_7090, n18_adj_7091, n24_adj_7092, 
        n18_adj_7093, n4_adj_7094, n20_adj_7095, n3_adj_7096, n26_adj_7097, 
        n22_adj_7098, n21_adj_7099, n18_adj_7100, n24_adj_7101, n18_adj_7102, 
        n4_adj_7103, n16_adj_7104, n17_adj_7105, n20_adj_7106, n5_adj_7107, 
        n3_adj_7108, n26_adj_7109, n22_adj_7110, n21_adj_7111, n18_adj_7112, 
        n24_adj_7113, n18_adj_7114, n4_adj_7115, n16_adj_7116, n17_adj_7117, 
        n20_adj_7118, n5_adj_7119, n3_adj_7120, n26_adj_7121, n22_adj_7122, 
        n21_adj_7123, n18_adj_7124, n24_adj_7125, n18_adj_7126, n4_adj_7127, 
        n16_adj_7128, n17_adj_7129, n20_adj_7130, n5_adj_7131, n3_adj_7132, 
        n26_adj_7133, n22_adj_7134, n21_adj_7135, n18_adj_7136, n24_adj_7137, 
        n18_adj_7138, n4_adj_7139, n16_adj_7140, n17_adj_7141, n20_adj_7142, 
        n5_adj_7143, n3_adj_7144, n26_adj_7145, n24_adj_7146, n18_adj_7147, 
        n4_adj_7148, n20_adj_7149;
    
    LUT4 i13_4_lut (.A(n3_c), .B(n26), .C(n22), .D(n21_c), .Z(\spi_data_out_r[26] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 Select_4060_i3_2_lut (.A(\spi_data_out_r_39__N_1168[26] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_c)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4060_i3_2_lut.init = 16'h8888;
    FD1P3IX mode__i0 (.D(n29762), .SP(clk_enable_288), .CD(n29239), .CK(clk), 
            .Q(mode_adj_181[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i0.GSR = "DISABLED";
    LUT4 i12_4_lut (.A(n18), .B(n24), .C(n18_adj_6759), .D(n4_c), .Z(n26)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 Select_4071_i5_2_lut (.A(\spi_data_out_r_39__N_1636[15] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4071_i5_2_lut.init = 16'h8888;
    LUT4 i8_4_lut (.A(\spi_data_out_r_39__N_4835[26] ), .B(n16), .C(n17_c), 
         .D(spi_data_out_r_39__N_4875), .Z(n22)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut.init = 16'hfefc;
    LUT4 Select_4060_i21_2_lut (.A(\spi_data_out_r_39__N_5513[26] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_c)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4060_i21_2_lut.init = 16'h8888;
    LUT4 Select_4060_i18_2_lut (.A(\spi_data_out_r_39__N_4496[26] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4060_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut (.A(\spi_data_out_r_39__N_3818[26] ), .B(n20_c), .C(n5_adj_6760), 
         .D(spi_data_out_r_39__N_3858), .Z(n24)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut.init = 16'hfefc;
    LUT4 i4_4_lut (.A(\spi_data_out_r_39__N_2104[26] ), .B(\spi_data_out_r_39__N_1870[26] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6759)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut.init = 16'heca0;
    LUT4 Select_4060_i4_2_lut (.A(\spi_data_out_r_39__N_1402[26] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_c)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4060_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut (.A(\spi_data_out_r_39__N_2338[26] ), .B(\spi_data_out_r_39__N_5174[26] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut.init = 16'heca0;
    LUT4 Select_4060_i5_2_lut (.A(\spi_data_out_r_39__N_1636[26] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6760)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4060_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut (.A(\spi_data_out_r_39__N_934[26] ), .B(spi_data_out_r_39__N_5852[26]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut.init = 16'heca0;
    LUT4 Select_4060_i17_2_lut (.A(\spi_data_out_r_39__N_4157[26] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_c)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4060_i17_2_lut.init = 16'h8888;
    LUT4 Select_4087_i1_2_lut_3_lut_4_lut (.A(mode_adj_181[2]), .B(mode_adj_181[1]), 
         .C(pin_io_out_68), .D(mode_adj_181[0]), .Z(\quad_a[6] )) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam Select_4087_i1_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 RESET_N_6154_bdd_2_lut_3_lut (.A(mode_adj_181[2]), .B(mode_adj_181[1]), 
         .C(mode_adj_181[0]), .Z(n28811)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam RESET_N_6154_bdd_2_lut_3_lut.init = 16'hbfbf;
    LUT4 i13_4_lut_adj_573 (.A(n3_adj_6761), .B(n26_adj_6762), .C(n22_adj_6763), 
         .D(n21_adj_6764), .Z(\spi_data_out_r[27] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_573.init = 16'hfffe;
    LUT4 Select_4094_i1_2_lut_3_lut_4_lut (.A(mode_adj_181[2]), .B(mode_adj_181[1]), 
         .C(pin_io_out_69), .D(mode_adj_181[0]), .Z(\quad_b[6] )) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam Select_4094_i1_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 Select_4059_i3_2_lut (.A(\spi_data_out_r_39__N_1168[27] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_6761)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4059_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_574 (.A(n18_adj_6765), .B(n24_adj_6766), .C(n18_adj_6767), 
         .D(n4_adj_6768), .Z(n26_adj_6762)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_574.init = 16'hfffe;
    LUT4 i8_4_lut_adj_575 (.A(\spi_data_out_r_39__N_4835[27] ), .B(n16_adj_6769), 
         .C(n17_adj_6770), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6763)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_575.init = 16'hfefc;
    LUT4 Select_4059_i21_2_lut (.A(\spi_data_out_r_39__N_5513[27] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6764)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4059_i21_2_lut.init = 16'h8888;
    LUT4 i8_4_lut_adj_576 (.A(\spi_data_out_r_39__N_4835[21] ), .B(n16_adj_6771), 
         .C(n17_adj_6772), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6773)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_576.init = 16'hfefc;
    LUT4 Select_4059_i18_2_lut (.A(\spi_data_out_r_39__N_4496[27] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6765)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4059_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_577 (.A(\spi_data_out_r_39__N_3818[27] ), .B(n20_adj_6774), 
         .C(n5_adj_6775), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_6766)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_577.init = 16'hfefc;
    LUT4 i4_4_lut_adj_578 (.A(\spi_data_out_r_39__N_2104[27] ), .B(\spi_data_out_r_39__N_1870[27] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6767)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_578.init = 16'heca0;
    LUT4 Select_4059_i4_2_lut (.A(\spi_data_out_r_39__N_1402[27] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6768)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4059_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_579 (.A(\spi_data_out_r_39__N_2338[27] ), .B(\spi_data_out_r_39__N_5174[27] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_6774)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_579.init = 16'heca0;
    LUT4 Select_4059_i5_2_lut (.A(\spi_data_out_r_39__N_1636[27] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6775)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4059_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_580 (.A(\spi_data_out_r_39__N_934[27] ), .B(spi_data_out_r_39__N_5852[27]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6769)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_580.init = 16'heca0;
    LUT4 Select_4059_i17_2_lut (.A(\spi_data_out_r_39__N_4157[27] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6770)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4059_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_581 (.A(n3_adj_6776), .B(n26_adj_6777), .C(n22_adj_6778), 
         .D(n21_adj_6779), .Z(\spi_data_out_r[28] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_581.init = 16'hfffe;
    LUT4 Select_4058_i3_2_lut (.A(\spi_data_out_r_39__N_1168[28] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_6776)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4058_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_582 (.A(n18_adj_6780), .B(n24_adj_6781), .C(n18_adj_6782), 
         .D(n4_adj_6783), .Z(n26_adj_6777)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_582.init = 16'hfffe;
    FD1S3AX SLO_buf_i1 (.D(SLO[0]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i1.GSR = "DISABLED";
    FD1P3AX SLO_i0 (.D(pin_io_out_68), .SP(clk_1MHz_derived_322_enable_20), 
            .CK(clk_1MHz_derived_322), .Q(SLO[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i0 (.D(\spi_data_out_r_39__N_6114[0] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_5852[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i0.GSR = "DISABLED";
    LUT4 i8_4_lut_adj_583 (.A(\spi_data_out_r_39__N_4835[28] ), .B(n16_adj_6784), 
         .C(n17_adj_6785), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6778)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_583.init = 16'hfefc;
    FD1P3IX Cnt_NSL__i0 (.D(n1290[0]), .SP(clk_1MHz_enable_367), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i0.GSR = "DISABLED";
    FD1P3IX Cnt__i0 (.D(n199[0]), .SP(clk_1MHz_enable_374), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i0.GSR = "DISABLED";
    LUT4 Select_4058_i21_2_lut (.A(\spi_data_out_r_39__N_5513[28] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6779)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4058_i21_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_584 (.A(\spi_data_out_r_39__N_934[15] ), .B(spi_data_out_r_39__N_5852[15]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6786)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_584.init = 16'heca0;
    LUT4 Select_4071_i17_2_lut (.A(\spi_data_out_r_39__N_4157[15] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6787)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4071_i17_2_lut.init = 16'h8888;
    LUT4 Select_4058_i18_2_lut (.A(\spi_data_out_r_39__N_4496[28] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6780)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4058_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_585 (.A(\spi_data_out_r_39__N_3818[28] ), .B(n20_adj_6788), 
         .C(n5_adj_6789), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_6781)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_585.init = 16'hfefc;
    LUT4 i4_4_lut_adj_586 (.A(\spi_data_out_r_39__N_2104[28] ), .B(\spi_data_out_r_39__N_1870[28] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6782)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_586.init = 16'heca0;
    LUT4 Select_4058_i4_2_lut (.A(\spi_data_out_r_39__N_1402[28] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6783)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4058_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_587 (.A(\spi_data_out_r_39__N_2338[28] ), .B(\spi_data_out_r_39__N_5174[28] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_6788)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_587.init = 16'heca0;
    LUT4 Select_4065_i5_2_lut (.A(\spi_data_out_r_39__N_1636[21] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6790)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4065_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_588 (.A(\spi_data_out_r_39__N_934[21] ), .B(spi_data_out_r_39__N_5852[21]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6771)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_588.init = 16'heca0;
    LUT4 Select_4065_i17_2_lut (.A(\spi_data_out_r_39__N_4157[21] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6772)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4065_i17_2_lut.init = 16'h8888;
    LUT4 Select_4058_i5_2_lut (.A(\spi_data_out_r_39__N_1636[28] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6789)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4058_i5_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_589 (.A(n3_adj_6791), .B(n26_adj_6792), .C(n22_adj_6793), 
         .D(n21_adj_6794), .Z(\spi_data_out_r[22] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_589.init = 16'hfffe;
    LUT4 Select_4064_i3_2_lut (.A(\spi_data_out_r_39__N_1168[22] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_6791)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4064_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_590 (.A(n18_adj_6795), .B(n24_adj_6796), .C(n18_adj_6797), 
         .D(n4_adj_6798), .Z(n26_adj_6792)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_590.init = 16'hfffe;
    LUT4 i8_4_lut_adj_591 (.A(\spi_data_out_r_39__N_4835[22] ), .B(n16_adj_6799), 
         .C(n17_adj_6800), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6793)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_591.init = 16'hfefc;
    LUT4 Select_4064_i21_2_lut (.A(\spi_data_out_r_39__N_5513[22] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6794)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4064_i21_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_592 (.A(\spi_data_out_r_39__N_934[28] ), .B(spi_data_out_r_39__N_5852[28]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6784)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_592.init = 16'heca0;
    LUT4 Select_4058_i17_2_lut (.A(\spi_data_out_r_39__N_4157[28] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6785)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4058_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_593 (.A(n3_adj_6801), .B(n26_adj_6802), .C(n22_adj_6803), 
         .D(n21_adj_6804), .Z(\spi_data_out_r[29] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_593.init = 16'hfffe;
    LUT4 Select_4064_i18_2_lut (.A(\spi_data_out_r_39__N_4496[22] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6795)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4064_i18_2_lut.init = 16'h8888;
    LUT4 Select_4057_i3_2_lut (.A(\spi_data_out_r_39__N_1168[29] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_6801)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4057_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_594 (.A(n18_adj_6805), .B(n24_adj_6806), .C(n18_adj_6807), 
         .D(n4_adj_6808), .Z(n26_adj_6802)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_594.init = 16'hfffe;
    LUT4 i8_4_lut_adj_595 (.A(\spi_data_out_r_39__N_4835[29] ), .B(n16_adj_6809), 
         .C(n17_adj_6810), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6803)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_595.init = 16'hfefc;
    LUT4 Select_4057_i21_2_lut (.A(\spi_data_out_r_39__N_5513[29] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6804)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4057_i21_2_lut.init = 16'h8888;
    LUT4 Select_4057_i18_2_lut (.A(\spi_data_out_r_39__N_4496[29] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6805)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4057_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_596 (.A(\spi_data_out_r_39__N_3818[29] ), .B(n20_adj_6811), 
         .C(n5_adj_6812), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_6806)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_596.init = 16'hfefc;
    LUT4 i10_4_lut_adj_597 (.A(\spi_data_out_r_39__N_3818[22] ), .B(n20_adj_6813), 
         .C(n5_adj_6814), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_6796)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_597.init = 16'hfefc;
    PFUMX i23073 (.BLUT(n28796), .ALUT(n28795), .C0(n19545), .Z(n28797));
    LUT4 i4_4_lut_adj_598 (.A(\spi_data_out_r_39__N_2104[29] ), .B(\spi_data_out_r_39__N_1870[29] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6807)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_598.init = 16'heca0;
    LUT4 i4_4_lut_adj_599 (.A(\spi_data_out_r_39__N_2104[22] ), .B(\spi_data_out_r_39__N_1870[22] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6797)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_599.init = 16'heca0;
    LUT4 Select_4064_i4_2_lut (.A(\spi_data_out_r_39__N_1402[22] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6798)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4064_i4_2_lut.init = 16'h8888;
    LUT4 Select_4057_i4_2_lut (.A(\spi_data_out_r_39__N_1402[29] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6808)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4057_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_600 (.A(\spi_data_out_r_39__N_2338[29] ), .B(\spi_data_out_r_39__N_5174[29] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_6811)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_600.init = 16'heca0;
    LUT4 Select_4057_i5_2_lut (.A(\spi_data_out_r_39__N_1636[29] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6812)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4057_i5_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_601 (.A(\spi_data_out_r_39__N_2338[22] ), .B(\spi_data_out_r_39__N_5174[22] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_6813)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_601.init = 16'heca0;
    LUT4 i2_4_lut_adj_602 (.A(\spi_data_out_r_39__N_934[29] ), .B(spi_data_out_r_39__N_5852[29]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6809)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_602.init = 16'heca0;
    FD1S3IX i159_483 (.D(n29087), .CK(clk), .CD(n29239), .Q(spi_data_out_r_39__N_5892)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam i159_483.GSR = "DISABLED";
    LUT4 Select_4057_i17_2_lut (.A(\spi_data_out_r_39__N_4157[29] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6810)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4057_i17_2_lut.init = 16'h8888;
    LUT4 Select_4064_i5_2_lut (.A(\spi_data_out_r_39__N_1636[22] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6814)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4064_i5_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_603 (.A(n3_adj_6815), .B(n26_adj_6816), .C(n22_adj_6817), 
         .D(n21_adj_6818), .Z(\spi_data_out_r[30] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_603.init = 16'hfffe;
    LUT4 Select_4056_i3_2_lut (.A(\spi_data_out_r_39__N_1168[30] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_6815)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4056_i3_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_604 (.A(\spi_data_out_r_39__N_934[22] ), .B(spi_data_out_r_39__N_5852[22]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6799)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_604.init = 16'heca0;
    LUT4 i12_4_lut_adj_605 (.A(n18_adj_6819), .B(n24_adj_6820), .C(n18_adj_6821), 
         .D(n4_adj_6822), .Z(n26_adj_6816)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_605.init = 16'hfffe;
    LUT4 i8_4_lut_adj_606 (.A(\spi_data_out_r_39__N_4835[30] ), .B(n16_adj_6823), 
         .C(n17_adj_6824), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6817)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_606.init = 16'hfefc;
    LUT4 Select_4056_i21_2_lut (.A(\spi_data_out_r_39__N_5513[30] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6818)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4056_i21_2_lut.init = 16'h8888;
    LUT4 Select_4064_i17_2_lut (.A(\spi_data_out_r_39__N_4157[22] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6800)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4064_i17_2_lut.init = 16'h8888;
    LUT4 Select_4056_i18_2_lut (.A(\spi_data_out_r_39__N_4496[30] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6819)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4056_i18_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_607 (.A(n3_adj_6825), .B(n26_adj_6826), .C(n22_adj_6827), 
         .D(n21_adj_6828), .Z(\spi_data_out_r[23] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_607.init = 16'hfffe;
    LUT4 i10_4_lut_adj_608 (.A(\spi_data_out_r_39__N_3818[30] ), .B(n20_adj_6829), 
         .C(n5_adj_6830), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_6820)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_608.init = 16'hfefc;
    FD1P3IX digital_output_r_481 (.D(\spi_data_r[0] ), .SP(clk_enable_198), 
            .CD(n29239), .CK(clk), .Q(digital_output_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam digital_output_r_481.GSR = "DISABLED";
    LUT4 Select_4063_i3_2_lut (.A(\spi_data_out_r_39__N_1168[23] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_6825)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4063_i3_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_609 (.A(\spi_data_out_r_39__N_2104[30] ), .B(\spi_data_out_r_39__N_1870[30] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6821)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_609.init = 16'heca0;
    LUT4 i12_4_lut_adj_610 (.A(n18_adj_6831), .B(n24_adj_6832), .C(n18_adj_6833), 
         .D(n4_adj_6834), .Z(n26_adj_6826)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_610.init = 16'hfffe;
    LUT4 Select_4056_i4_2_lut (.A(\spi_data_out_r_39__N_1402[30] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6822)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4056_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_611 (.A(\spi_data_out_r_39__N_2338[30] ), .B(\spi_data_out_r_39__N_5174[30] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_6829)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_611.init = 16'heca0;
    LUT4 Select_4056_i5_2_lut (.A(\spi_data_out_r_39__N_1636[30] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6830)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4056_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_612 (.A(\spi_data_out_r_39__N_934[30] ), .B(spi_data_out_r_39__N_5852[30]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6823)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_612.init = 16'heca0;
    LUT4 Select_4056_i17_2_lut (.A(\spi_data_out_r_39__N_4157[30] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6824)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4056_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_613 (.A(n3_adj_6835), .B(n26_adj_6836), .C(n22_adj_6837), 
         .D(n21_adj_6838), .Z(\spi_data_out_r[31] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_613.init = 16'hfffe;
    LUT4 i8_4_lut_adj_614 (.A(\spi_data_out_r_39__N_4835[23] ), .B(n16_adj_6839), 
         .C(n17_adj_6840), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6827)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_614.init = 16'hfefc;
    LUT4 Select_4055_i3_2_lut (.A(\spi_data_out_r_39__N_1168[31] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_6835)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4055_i3_2_lut.init = 16'h8888;
    LUT4 Select_4063_i21_2_lut (.A(\spi_data_out_r_39__N_5513[23] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6828)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4063_i21_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_615 (.A(n3_adj_6841), .B(n26_adj_6842), .C(n22_adj_6843), 
         .D(n21_adj_6844), .Z(\spi_data_out_r[16] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_615.init = 16'hfffe;
    LUT4 Select_4070_i3_2_lut (.A(\spi_data_out_r_39__N_1168[16] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_6841)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4070_i3_2_lut.init = 16'h8888;
    LUT4 Select_4063_i18_2_lut (.A(\spi_data_out_r_39__N_4496[23] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6831)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4063_i18_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_616 (.A(n18_adj_6845), .B(n24_adj_6846), .C(n18_adj_6847), 
         .D(n4_adj_6848), .Z(n26_adj_6836)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_616.init = 16'hfffe;
    LUT4 i8_4_lut_adj_617 (.A(\spi_data_out_r_39__N_4835[31] ), .B(n16_adj_6849), 
         .C(n17_adj_6850), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6837)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_617.init = 16'hfefc;
    LUT4 i10_4_lut_adj_618 (.A(\spi_data_out_r_39__N_3818[23] ), .B(n20_adj_6851), 
         .C(n5_adj_6852), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_6832)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_618.init = 16'hfefc;
    LUT4 Select_4055_i21_2_lut (.A(\spi_data_out_r_39__N_5513[31] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6838)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4055_i21_2_lut.init = 16'h8888;
    LUT4 Select_4055_i18_2_lut (.A(\spi_data_out_r_39__N_4496[31] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6845)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4055_i18_2_lut.init = 16'h8888;
    LUT4 i22681_2_lut_rep_417 (.A(n19401), .B(resetn_c), .Z(clk_1MHz_enable_374)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i22681_2_lut_rep_417.init = 16'hbbbb;
    LUT4 i10_4_lut_adj_619 (.A(\spi_data_out_r_39__N_3818[31] ), .B(n20_adj_6853), 
         .C(n5_adj_6854), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_6846)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_619.init = 16'hfefc;
    LUT4 i22861_2_lut_2_lut_3_lut_4_lut (.A(n19401), .B(resetn_c), .C(n19545), 
         .D(n19439), .Z(clk_1MHz_enable_377)) /* synthesis lut_function=(!(A (C (D))+!A (B+(C (D))))) */ ;
    defparam i22861_2_lut_2_lut_3_lut_4_lut.init = 16'h0bbb;
    LUT4 i4_4_lut_adj_620 (.A(\spi_data_out_r_39__N_2104[31] ), .B(\spi_data_out_r_39__N_1870[31] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6847)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_620.init = 16'heca0;
    LUT4 Select_4055_i4_2_lut (.A(\spi_data_out_r_39__N_1402[31] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6848)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4055_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_621 (.A(\spi_data_out_r_39__N_2338[31] ), .B(\spi_data_out_r_39__N_5174[31] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_6853)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_621.init = 16'heca0;
    LUT4 Select_4055_i5_2_lut (.A(\spi_data_out_r_39__N_1636[31] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6854)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4055_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_622 (.A(\spi_data_out_r_39__N_934[31] ), .B(spi_data_out_r_39__N_5852[31]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6849)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_622.init = 16'heca0;
    LUT4 Select_4055_i17_2_lut (.A(\spi_data_out_r_39__N_4157[31] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6850)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4055_i17_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_623 (.A(\spi_data_out_r_39__N_4835[32] ), .B(n12), 
         .C(n8_c), .D(spi_data_out_r_39__N_4875), .Z(\spi_data_out_r[32] )) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_623.init = 16'hfefc;
    LUT4 i5_4_lut (.A(\spi_data_out_r_39__N_3818[32] ), .B(n10), .C(n21_adj_6855), 
         .D(spi_data_out_r_39__N_3858), .Z(n12)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut.init = 16'hfefc;
    LUT4 i1_4_lut (.A(spi_data_out_r_39__N_5852[32]), .B(\spi_data_out_r_39__N_5174[32] ), 
         .C(spi_data_out_r_39__N_5892), .D(spi_data_out_r_39__N_5214), .Z(n8_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut.init = 16'heca0;
    LUT4 i3_4_lut (.A(\spi_data_out_r_39__N_4496[32] ), .B(\spi_data_out_r_39__N_4157[32] ), 
         .C(spi_data_out_r_39__N_4536), .D(spi_data_out_r_39__N_4197), .Z(n10)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut.init = 16'heca0;
    LUT4 Select_4054_i21_2_lut (.A(\spi_data_out_r_39__N_5513[32] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6855)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4054_i21_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_624 (.A(\spi_data_out_r_39__N_4835[33] ), .B(n12_adj_6856), 
         .C(n8_adj_6857), .D(spi_data_out_r_39__N_4875), .Z(\spi_data_out_r[33] )) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_624.init = 16'hfefc;
    LUT4 i5_4_lut_adj_625 (.A(\spi_data_out_r_39__N_3818[33] ), .B(n10_adj_6858), 
         .C(n21_adj_6859), .D(spi_data_out_r_39__N_3858), .Z(n12_adj_6856)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_625.init = 16'hfefc;
    LUT4 i1_4_lut_adj_626 (.A(spi_data_out_r_39__N_5852[33]), .B(\spi_data_out_r_39__N_5174[33] ), 
         .C(spi_data_out_r_39__N_5892), .D(spi_data_out_r_39__N_5214), .Z(n8_adj_6857)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_626.init = 16'heca0;
    LUT4 i3_4_lut_adj_627 (.A(\spi_data_out_r_39__N_4496[33] ), .B(\spi_data_out_r_39__N_4157[33] ), 
         .C(spi_data_out_r_39__N_4536), .D(spi_data_out_r_39__N_4197), .Z(n10_adj_6858)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_627.init = 16'heca0;
    LUT4 Select_4053_i21_2_lut (.A(\spi_data_out_r_39__N_5513[33] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6859)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4053_i21_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_628 (.A(\spi_data_out_r_39__N_4835[34] ), .B(n12_adj_6860), 
         .C(n8_adj_6861), .D(spi_data_out_r_39__N_4875), .Z(\spi_data_out_r[34] )) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_628.init = 16'hfefc;
    LUT4 i5_4_lut_adj_629 (.A(\spi_data_out_r_39__N_3818[34] ), .B(n10_adj_6862), 
         .C(n21_adj_6863), .D(spi_data_out_r_39__N_3858), .Z(n12_adj_6860)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_629.init = 16'hfefc;
    LUT4 i1_4_lut_adj_630 (.A(spi_data_out_r_39__N_5852[34]), .B(\spi_data_out_r_39__N_5174[34] ), 
         .C(spi_data_out_r_39__N_5892), .D(spi_data_out_r_39__N_5214), .Z(n8_adj_6861)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_630.init = 16'heca0;
    LUT4 i3_4_lut_adj_631 (.A(\spi_data_out_r_39__N_4496[34] ), .B(\spi_data_out_r_39__N_4157[34] ), 
         .C(spi_data_out_r_39__N_4536), .D(spi_data_out_r_39__N_4197), .Z(n10_adj_6862)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_631.init = 16'heca0;
    LUT4 i4_4_lut_adj_632 (.A(\spi_data_out_r_39__N_2104[23] ), .B(\spi_data_out_r_39__N_1870[23] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6833)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_632.init = 16'heca0;
    LUT4 Select_4052_i21_2_lut (.A(\spi_data_out_r_39__N_5513[34] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6863)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4052_i21_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_633 (.A(\spi_data_out_r_39__N_4835[35] ), .B(n12_adj_6864), 
         .C(n8_adj_6865), .D(spi_data_out_r_39__N_4875), .Z(\spi_data_out_r[35] )) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_633.init = 16'hfefc;
    LUT4 i5_4_lut_adj_634 (.A(\spi_data_out_r_39__N_3818[35] ), .B(n10_adj_6866), 
         .C(n21_adj_6867), .D(spi_data_out_r_39__N_3858), .Z(n12_adj_6864)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_634.init = 16'hfefc;
    LUT4 i1_4_lut_adj_635 (.A(spi_data_out_r_39__N_5852[35]), .B(\spi_data_out_r_39__N_5174[35] ), 
         .C(spi_data_out_r_39__N_5892), .D(spi_data_out_r_39__N_5214), .Z(n8_adj_6865)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_635.init = 16'heca0;
    LUT4 i3_4_lut_adj_636 (.A(\spi_data_out_r_39__N_4496[35] ), .B(\spi_data_out_r_39__N_4157[35] ), 
         .C(spi_data_out_r_39__N_4536), .D(spi_data_out_r_39__N_4197), .Z(n10_adj_6866)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_636.init = 16'heca0;
    LUT4 Select_4051_i21_2_lut (.A(\spi_data_out_r_39__N_5513[35] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6867)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4051_i21_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_637 (.A(\spi_data_out_r_39__N_4835[36] ), .B(n12_adj_6868), 
         .C(n8_adj_6869), .D(spi_data_out_r_39__N_4875), .Z(\spi_data_out_r[36] )) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_637.init = 16'hfefc;
    LUT4 i5_4_lut_adj_638 (.A(\spi_data_out_r_39__N_3818[36] ), .B(n10_adj_6870), 
         .C(n21_adj_6871), .D(spi_data_out_r_39__N_3858), .Z(n12_adj_6868)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_638.init = 16'hfefc;
    LUT4 i1_4_lut_adj_639 (.A(spi_data_out_r_39__N_5852[36]), .B(\spi_data_out_r_39__N_5174[36] ), 
         .C(spi_data_out_r_39__N_5892), .D(spi_data_out_r_39__N_5214), .Z(n8_adj_6869)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_639.init = 16'heca0;
    LUT4 i3_4_lut_adj_640 (.A(\spi_data_out_r_39__N_4496[36] ), .B(\spi_data_out_r_39__N_4157[36] ), 
         .C(spi_data_out_r_39__N_4536), .D(spi_data_out_r_39__N_4197), .Z(n10_adj_6870)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_640.init = 16'heca0;
    LUT4 Select_4050_i21_2_lut (.A(\spi_data_out_r_39__N_5513[36] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6871)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4050_i21_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_641 (.A(\spi_data_out_r_39__N_4835[37] ), .B(n12_adj_6872), 
         .C(n8_adj_6873), .D(spi_data_out_r_39__N_4875), .Z(\spi_data_out_r[37] )) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_641.init = 16'hfefc;
    LUT4 Select_4063_i4_2_lut (.A(\spi_data_out_r_39__N_1402[23] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6834)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4063_i4_2_lut.init = 16'h8888;
    LUT4 i5_4_lut_adj_642 (.A(\spi_data_out_r_39__N_3818[37] ), .B(n10_adj_6874), 
         .C(n21_adj_6875), .D(spi_data_out_r_39__N_3858), .Z(n12_adj_6872)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_642.init = 16'hfefc;
    LUT4 i1_4_lut_adj_643 (.A(spi_data_out_r_39__N_5852[37]), .B(\spi_data_out_r_39__N_5174[37] ), 
         .C(spi_data_out_r_39__N_5892), .D(spi_data_out_r_39__N_5214), .Z(n8_adj_6873)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_643.init = 16'heca0;
    LUT4 i3_4_lut_adj_644 (.A(\spi_data_out_r_39__N_4496[37] ), .B(\spi_data_out_r_39__N_4157[37] ), 
         .C(spi_data_out_r_39__N_4536), .D(spi_data_out_r_39__N_4197), .Z(n10_adj_6874)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_644.init = 16'heca0;
    LUT4 i6_4_lut_adj_645 (.A(\spi_data_out_r_39__N_2338[23] ), .B(\spi_data_out_r_39__N_5174[23] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_6851)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_645.init = 16'heca0;
    LUT4 Select_4049_i21_2_lut (.A(\spi_data_out_r_39__N_5513[37] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6875)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4049_i21_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_646 (.A(\spi_data_out_r_39__N_4835[38] ), .B(n12_adj_6876), 
         .C(n8_adj_6877), .D(spi_data_out_r_39__N_4875), .Z(\spi_data_out_r[38] )) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_646.init = 16'hfefc;
    LUT4 i5_4_lut_adj_647 (.A(\spi_data_out_r_39__N_3818[38] ), .B(n10_adj_6878), 
         .C(n21_adj_6879), .D(spi_data_out_r_39__N_3858), .Z(n12_adj_6876)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_647.init = 16'hfefc;
    LUT4 Select_4063_i5_2_lut (.A(\spi_data_out_r_39__N_1636[23] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6852)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4063_i5_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_648 (.A(spi_data_out_r_39__N_5852[38]), .B(\spi_data_out_r_39__N_5174[38] ), 
         .C(spi_data_out_r_39__N_5892), .D(spi_data_out_r_39__N_5214), .Z(n8_adj_6877)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_648.init = 16'heca0;
    LUT4 i3_4_lut_adj_649 (.A(\spi_data_out_r_39__N_4496[38] ), .B(\spi_data_out_r_39__N_4157[38] ), 
         .C(spi_data_out_r_39__N_4536), .D(spi_data_out_r_39__N_4197), .Z(n10_adj_6878)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_649.init = 16'heca0;
    LUT4 i2_4_lut_adj_650 (.A(\spi_data_out_r_39__N_934[23] ), .B(spi_data_out_r_39__N_5852[23]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6839)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_650.init = 16'heca0;
    LUT4 Select_4063_i17_2_lut (.A(\spi_data_out_r_39__N_4157[23] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6840)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4063_i17_2_lut.init = 16'h8888;
    LUT4 Select_4048_i21_2_lut (.A(\spi_data_out_r_39__N_5513[38] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6879)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4048_i21_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_651 (.A(\spi_data_out_r_39__N_4835[39] ), .B(n12_adj_6880), 
         .C(n8_adj_6881), .D(spi_data_out_r_39__N_4875), .Z(\spi_data_out_r[39] )) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i6_4_lut_adj_651.init = 16'hfefc;
    LUT4 i5_4_lut_adj_652 (.A(\spi_data_out_r_39__N_3818[39] ), .B(n10_adj_6882), 
         .C(n21_adj_6883), .D(spi_data_out_r_39__N_3858), .Z(n12_adj_6880)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i5_4_lut_adj_652.init = 16'hfefc;
    LUT4 i22933_2_lut_rep_543 (.A(Cnt[4]), .B(Cnt[1]), .Z(n29271)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i22933_2_lut_rep_543.init = 16'h7777;
    LUT4 i1_2_lut_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(n29192), .D(Cnt[5]), 
         .Z(n11795)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff7;
    LUT4 i1_4_lut_adj_653 (.A(spi_data_out_r_39__N_5852[39]), .B(\spi_data_out_r_39__N_5174[39] ), 
         .C(spi_data_out_r_39__N_5892), .D(spi_data_out_r_39__N_5214), .Z(n8_adj_6881)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_653.init = 16'heca0;
    LUT4 i3_4_lut_adj_654 (.A(\spi_data_out_r_39__N_4496[39] ), .B(\spi_data_out_r_39__N_4157[39] ), 
         .C(spi_data_out_r_39__N_4536), .D(spi_data_out_r_39__N_4197), .Z(n10_adj_6882)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_654.init = 16'heca0;
    LUT4 n19439_bdd_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(Cnt[5]), .D(MA_Temp), 
         .Z(n28796)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;
    defparam n19439_bdd_3_lut_4_lut.init = 16'hf708;
    LUT4 Select_4047_i21_2_lut (.A(\spi_data_out_r_39__N_5513[39] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6883)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4047_i21_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_655 (.A(n3_adj_6884), .B(n26_adj_6885), .C(n22_adj_6886), 
         .D(n21_adj_6887), .Z(\spi_data_out_r[24] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_655.init = 16'hfffe;
    LUT4 Select_4062_i3_2_lut (.A(\spi_data_out_r_39__N_1168[24] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_6884)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4062_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_656 (.A(n18_adj_6888), .B(n24_adj_6889), .C(n18_adj_6890), 
         .D(n4_adj_6891), .Z(n26_adj_6885)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_656.init = 16'hfffe;
    LUT4 i8_4_lut_adj_657 (.A(\spi_data_out_r_39__N_4835[24] ), .B(n16_adj_6892), 
         .C(n17_adj_6893), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6886)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_657.init = 16'hfefc;
    LUT4 Select_4062_i21_2_lut (.A(\spi_data_out_r_39__N_5513[24] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6887)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4062_i21_2_lut.init = 16'h8888;
    LUT4 Select_4062_i18_2_lut (.A(\spi_data_out_r_39__N_4496[24] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6888)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4062_i18_2_lut.init = 16'h8888;
    LUT4 i4775_3_lut_rep_425_4_lut (.A(mode_adj_181[0]), .B(n29267), .C(mode), 
         .D(n29191), .Z(n29153)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;
    defparam i4775_3_lut_rep_425_4_lut.init = 16'h00fb;
    LUT4 i10_4_lut_adj_658 (.A(\spi_data_out_r_39__N_3818[24] ), .B(n20_adj_6894), 
         .C(n5_adj_6895), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_6889)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_658.init = 16'hfefc;
    LUT4 i1_2_lut_rep_547 (.A(Cnt[6]), .B(Cnt[7]), .Z(n29275)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_547.init = 16'heeee;
    LUT4 i2_3_lut_rep_464_4_lut (.A(Cnt[6]), .B(Cnt[7]), .C(Cnt[0]), .D(n27387), 
         .Z(n29192)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_464_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_428_4_lut (.A(n27387), .B(Cnt[0]), .C(n29275), .D(Cnt[5]), 
         .Z(n29156)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_rep_428_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_549 (.A(mode_adj_181[1]), .B(mode_adj_181[2]), .Z(n29277)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_rep_549.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_467_3_lut (.A(mode_adj_181[1]), .B(mode_adj_181[2]), 
         .C(mode_adj_181[0]), .Z(n29195)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_rep_467_3_lut.init = 16'hbfbf;
    LUT4 equal_163_i6_1_lut_2_lut_3_lut (.A(mode_adj_181[1]), .B(mode_adj_181[2]), 
         .C(mode_adj_181[0]), .Z(MA_Temp_N_5983)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam equal_163_i6_1_lut_2_lut_3_lut.init = 16'h4040;
    LUT4 i4_4_lut_adj_659 (.A(\spi_data_out_r_39__N_2104[24] ), .B(\spi_data_out_r_39__N_1870[24] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6890)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_659.init = 16'heca0;
    LUT4 Select_3870_i7_3_lut_4_lut (.A(mode_adj_181[0]), .B(n29277), .C(n29293), 
         .D(\cs_decoded[12] ), .Z(n8652)) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam Select_3870_i7_3_lut_4_lut.init = 16'hf222;
    LUT4 i1_2_lut_3_lut (.A(mode_adj_181[1]), .B(mode_adj_181[2]), .C(mode_adj_181[0]), 
         .Z(n13378)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_3_lut.init = 16'hfbfb;
    LUT4 Select_3850_i1_2_lut_3_lut_4_lut (.A(mode_adj_181[1]), .B(mode_adj_181[2]), 
         .C(NSL), .D(mode_adj_181[0]), .Z(n1)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam Select_3850_i1_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i4826_2_lut_3_lut_4_lut (.A(mode_adj_181[1]), .B(mode_adj_181[2]), 
         .C(clk_1MHz_derived_322_enable_46), .D(mode_adj_181[0]), .Z(clk_1MHz_derived_322_enable_20)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i4826_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i22770_2_lut_3_lut_3_lut_4_lut (.A(mode_adj_181[1]), .B(mode_adj_181[2]), 
         .C(mode_adj_181[0]), .D(n29293), .Z(n8651)) /* synthesis lut_function=(!(A (D)+!A (B (C+(D))+!B (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i22770_2_lut_3_lut_3_lut_4_lut.init = 16'h00bf;
    LUT4 i22675_2_lut_rep_550 (.A(MA_Temp), .B(clk_1MHz), .Z(clk_1MHz_derived_322)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[13:34])
    defparam i22675_2_lut_rep_550.init = 16'h7777;
    LUT4 Select_3847_i1_2_lut_3_lut (.A(MA_Temp), .B(clk_1MHz), .C(mode_adj_181[2]), 
         .Z(n1_adj_171)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[13:34])
    defparam Select_3847_i1_2_lut_3_lut.init = 16'h7070;
    LUT4 Select_4065_i21_2_lut (.A(\spi_data_out_r_39__N_5513[21] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6897)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4065_i21_2_lut.init = 16'h8888;
    LUT4 Select_4062_i4_2_lut (.A(\spi_data_out_r_39__N_1402[24] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6891)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4062_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_660 (.A(\spi_data_out_r_39__N_2338[24] ), .B(\spi_data_out_r_39__N_5174[24] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_6894)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_660.init = 16'heca0;
    LUT4 Select_4062_i5_2_lut (.A(\spi_data_out_r_39__N_1636[24] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6895)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4062_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_661 (.A(\spi_data_out_r_39__N_934[24] ), .B(spi_data_out_r_39__N_5852[24]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6892)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_661.init = 16'heca0;
    LUT4 Select_4062_i17_2_lut (.A(\spi_data_out_r_39__N_4157[24] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6893)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4062_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_662 (.A(n3_adj_6898), .B(n26_adj_6899), .C(n22_adj_6900), 
         .D(n21_adj_6901), .Z(\spi_data_out_r[25] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_662.init = 16'hfffe;
    LUT4 Select_4061_i3_2_lut (.A(\spi_data_out_r_39__N_1168[25] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_6898)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4061_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_663 (.A(n18_adj_6902), .B(n24_adj_6903), .C(n18_adj_6904), 
         .D(n4_adj_6905), .Z(n26_adj_6899)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_663.init = 16'hfffe;
    LUT4 i8_4_lut_adj_664 (.A(\spi_data_out_r_39__N_4835[25] ), .B(n16_adj_6906), 
         .C(n17_adj_6907), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6900)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_664.init = 16'hfefc;
    LUT4 Select_4061_i21_2_lut (.A(\spi_data_out_r_39__N_5513[25] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6901)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4061_i21_2_lut.init = 16'h8888;
    LUT4 Select_4061_i18_2_lut (.A(\spi_data_out_r_39__N_4496[25] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6902)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4061_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_665 (.A(\spi_data_out_r_39__N_3818[25] ), .B(n20_adj_6908), 
         .C(n5_adj_6909), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_6903)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_665.init = 16'hfefc;
    LUT4 i4_4_lut_adj_666 (.A(\spi_data_out_r_39__N_2104[25] ), .B(\spi_data_out_r_39__N_1870[25] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6904)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_666.init = 16'heca0;
    LUT4 Select_4061_i4_2_lut (.A(\spi_data_out_r_39__N_1402[25] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6905)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4061_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_667 (.A(\spi_data_out_r_39__N_2338[25] ), .B(\spi_data_out_r_39__N_5174[25] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_6908)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_667.init = 16'heca0;
    CCU2D add_551_13 (.A0(Cnt_NSL[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25044), 
          .S0(n1290[11]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_13.INIT0 = 16'h5aaa;
    defparam add_551_13.INIT1 = 16'h0000;
    defparam add_551_13.INJECT1_0 = "NO";
    defparam add_551_13.INJECT1_1 = "NO";
    CCU2D add_551_11 (.A0(Cnt_NSL[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25043), .COUT(n25044), .S0(n1290[9]), .S1(n1290[10]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_11.INIT0 = 16'h5aaa;
    defparam add_551_11.INIT1 = 16'h5aaa;
    defparam add_551_11.INJECT1_0 = "NO";
    defparam add_551_11.INJECT1_1 = "NO";
    CCU2D add_551_9 (.A0(Cnt_NSL[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25042), .COUT(n25043), .S0(n1290[7]), .S1(n1290[8]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_9.INIT0 = 16'h5aaa;
    defparam add_551_9.INIT1 = 16'h5aaa;
    defparam add_551_9.INJECT1_0 = "NO";
    defparam add_551_9.INJECT1_1 = "NO";
    LUT4 i117_4_lut (.A(n29156), .B(n13378), .C(Cnt[1]), .D(Cnt[4]), 
         .Z(clk_1MHz_derived_322_enable_46)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(132[15:49])
    defparam i117_4_lut.init = 16'h3332;
    LUT4 Select_4061_i5_2_lut (.A(\spi_data_out_r_39__N_1636[25] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6909)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4061_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_668 (.A(\spi_data_out_r_39__N_934[25] ), .B(spi_data_out_r_39__N_5852[25]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6906)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_668.init = 16'heca0;
    CCU2D add_551_7 (.A0(Cnt_NSL[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25041), .COUT(n25042), .S0(n1290[5]), .S1(n1290[6]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_7.INIT0 = 16'h5aaa;
    defparam add_551_7.INIT1 = 16'h5aaa;
    defparam add_551_7.INJECT1_0 = "NO";
    defparam add_551_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut (.A(Cnt[2]), .B(Cnt[3]), .Z(n27387)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 Select_4061_i17_2_lut (.A(\spi_data_out_r_39__N_4157[25] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6907)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4061_i17_2_lut.init = 16'h8888;
    CCU2D add_551_5 (.A0(Cnt_NSL[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25040), .COUT(n25041), .S0(n1290[3]), .S1(n1290[4]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_5.INIT0 = 16'h5aaa;
    defparam add_551_5.INIT1 = 16'h5aaa;
    defparam add_551_5.INJECT1_0 = "NO";
    defparam add_551_5.INJECT1_1 = "NO";
    FD1P3AX NSL_476 (.D(NSL_N_6180), .SP(clk_1MHz_enable_247), .CK(clk_1MHz), 
            .Q(NSL)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam NSL_476.GSR = "DISABLED";
    CCU2D add_551_3 (.A0(Cnt_NSL[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25039), .COUT(n25040), .S0(n1290[1]), .S1(n1290[2]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_3.INIT0 = 16'h5aaa;
    defparam add_551_3.INIT1 = 16'h5aaa;
    defparam add_551_3.INJECT1_0 = "NO";
    defparam add_551_3.INJECT1_1 = "NO";
    LUT4 i14475_3_lut (.A(n19545), .B(resetn_c), .C(n19401), .Z(clk_1MHz_enable_247)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B))) */ ;
    defparam i14475_3_lut.init = 16'h4c4c;
    LUT4 i22672_4_lut (.A(NSL), .B(n19401), .C(n19545), .D(n11795), 
         .Z(NSL_N_6180)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C+(D))))) */ ;
    defparam i22672_4_lut.init = 16'h3b37;
    CCU2D add_551_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n25039), .S1(n1290[0]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_1.INIT0 = 16'hF000;
    defparam add_551_1.INIT1 = 16'h5555;
    defparam add_551_1.INJECT1_0 = "NO";
    defparam add_551_1.INJECT1_1 = "NO";
    FD1P3IX mode__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_288), .CD(n29239), 
            .CK(clk), .Q(mode_adj_181[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i2.GSR = "DISABLED";
    FD1P3IX mode__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_288), .CD(n29239), 
            .CK(clk), .Q(mode_adj_181[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i1.GSR = "DISABLED";
    CCU2D add_552_9 (.A0(Cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25038), 
          .S0(n153[7]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_9.INIT0 = 16'h5aaa;
    defparam add_552_9.INIT1 = 16'h0000;
    defparam add_552_9.INJECT1_0 = "NO";
    defparam add_552_9.INJECT1_1 = "NO";
    LUT4 i12_4_lut_adj_669 (.A(n18_adj_6910), .B(n24_adj_6911), .C(n18_adj_6912), 
         .D(n4_adj_6913), .Z(n26_adj_6842)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_669.init = 16'hfffe;
    LUT4 i8_4_lut_adj_670 (.A(\spi_data_out_r_39__N_4835[16] ), .B(n16_adj_6914), 
         .C(n17_adj_6915), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6843)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_670.init = 16'hfefc;
    LUT4 Select_4084_i13_2_lut (.A(\spi_data_out_r_39__N_2856[2] ), .B(clear_intrpt), 
         .Z(n13)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4084_i13_2_lut.init = 16'h8888;
    LUT4 Select_4084_i4_2_lut (.A(\spi_data_out_r_39__N_1402[2] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4084_i4_2_lut.init = 16'h8888;
    FD1S3AX SLO_buf_i2 (.D(SLO[1]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i2.GSR = "DISABLED";
    FD1S3AX SLO_buf_i3 (.D(SLO[2]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i3.GSR = "DISABLED";
    FD1S3AX SLO_buf_i4 (.D(SLO[3]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i4.GSR = "DISABLED";
    FD1S3AX SLO_buf_i5 (.D(SLO[4]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i5.GSR = "DISABLED";
    FD1S3AX SLO_buf_i6 (.D(SLO[5]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i6.GSR = "DISABLED";
    FD1S3AX SLO_buf_i7 (.D(SLO[6]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i7.GSR = "DISABLED";
    FD1S3AX SLO_buf_i8 (.D(SLO[7]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i8.GSR = "DISABLED";
    FD1S3AX SLO_buf_i9 (.D(SLO[8]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i9.GSR = "DISABLED";
    FD1S3AX SLO_buf_i10 (.D(SLO[9]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i10.GSR = "DISABLED";
    FD1S3AX SLO_buf_i11 (.D(SLO[10]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i11.GSR = "DISABLED";
    FD1S3AX SLO_buf_i12 (.D(SLO[11]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i12.GSR = "DISABLED";
    FD1S3AX SLO_buf_i13 (.D(SLO[12]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i13.GSR = "DISABLED";
    FD1S3AX SLO_buf_i14 (.D(SLO[13]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i14.GSR = "DISABLED";
    FD1S3AX SLO_buf_i15 (.D(SLO[14]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i15.GSR = "DISABLED";
    FD1S3AX SLO_buf_i16 (.D(SLO[15]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i16.GSR = "DISABLED";
    FD1S3AX SLO_buf_i17 (.D(SLO[16]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i17.GSR = "DISABLED";
    FD1S3AX SLO_buf_i18 (.D(SLO[17]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i18.GSR = "DISABLED";
    FD1S3AX SLO_buf_i19 (.D(SLO[18]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i19.GSR = "DISABLED";
    FD1S3AX SLO_buf_i20 (.D(SLO[19]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i20.GSR = "DISABLED";
    FD1S3AX SLO_buf_i21 (.D(SLO[20]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i21.GSR = "DISABLED";
    FD1S3AX SLO_buf_i22 (.D(SLO[21]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i22.GSR = "DISABLED";
    FD1S3AX SLO_buf_i23 (.D(SLO[22]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i23.GSR = "DISABLED";
    FD1S3AX SLO_buf_i24 (.D(SLO[23]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i24.GSR = "DISABLED";
    FD1S3AX SLO_buf_i25 (.D(SLO[24]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i25.GSR = "DISABLED";
    FD1S3AX SLO_buf_i26 (.D(SLO[25]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i26.GSR = "DISABLED";
    FD1S3AX SLO_buf_i27 (.D(SLO[26]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i27.GSR = "DISABLED";
    FD1S3AX SLO_buf_i28 (.D(SLO[27]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i28.GSR = "DISABLED";
    FD1S3AX SLO_buf_i29 (.D(SLO[28]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i29.GSR = "DISABLED";
    FD1S3AX SLO_buf_i30 (.D(SLO[29]), .CK(MA_Temp_N_5969), .Q(\SLO_buf[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i30.GSR = "DISABLED";
    FD1S3AX SLO_buf_i31 (.D(SLO[30]), .CK(MA_Temp_N_5969), .Q(SLO_buf[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i31.GSR = "DISABLED";
    FD1S3AX SLO_buf_i32 (.D(SLO[31]), .CK(MA_Temp_N_5969), .Q(SLO_buf[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i32.GSR = "DISABLED";
    FD1S3AX SLO_buf_i33 (.D(SLO[32]), .CK(MA_Temp_N_5969), .Q(SLO_buf[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i33.GSR = "DISABLED";
    FD1S3AX SLO_buf_i34 (.D(SLO[33]), .CK(MA_Temp_N_5969), .Q(SLO_buf[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i34.GSR = "DISABLED";
    FD1S3AX SLO_buf_i35 (.D(SLO[34]), .CK(MA_Temp_N_5969), .Q(SLO_buf[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i35.GSR = "DISABLED";
    FD1S3AX SLO_buf_i36 (.D(SLO[35]), .CK(MA_Temp_N_5969), .Q(SLO_buf[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i36.GSR = "DISABLED";
    FD1S3AX SLO_buf_i37 (.D(SLO[36]), .CK(MA_Temp_N_5969), .Q(SLO_buf[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i37.GSR = "DISABLED";
    FD1S3AX SLO_buf_i38 (.D(SLO[37]), .CK(MA_Temp_N_5969), .Q(SLO_buf[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i38.GSR = "DISABLED";
    FD1S3AX SLO_buf_i39 (.D(SLO[38]), .CK(MA_Temp_N_5969), .Q(SLO_buf[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i39.GSR = "DISABLED";
    FD1S3AX SLO_buf_i40 (.D(SLO[39]), .CK(MA_Temp_N_5969), .Q(SLO_buf[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i40.GSR = "DISABLED";
    FD1S3AX SLO_buf_i41 (.D(SLO[40]), .CK(MA_Temp_N_5969), .Q(SLO_buf[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i41.GSR = "DISABLED";
    FD1S3AX SLO_buf_i42 (.D(SLO[41]), .CK(MA_Temp_N_5969), .Q(SLO_buf[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i42.GSR = "DISABLED";
    FD1S3AX SLO_buf_i43 (.D(SLO[42]), .CK(MA_Temp_N_5969), .Q(SLO_buf[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i43.GSR = "DISABLED";
    FD1S3AX SLO_buf_i44 (.D(SLO[43]), .CK(MA_Temp_N_5969), .Q(SLO_buf[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i44.GSR = "DISABLED";
    FD1S3AX SLO_buf_i45 (.D(SLO[44]), .CK(MA_Temp_N_5969), .Q(SLO_buf[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i45.GSR = "DISABLED";
    FD1S3AX SLO_buf_i46 (.D(SLO[45]), .CK(MA_Temp_N_5969), .Q(SLO_buf[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i46.GSR = "DISABLED";
    FD1P3AX SLO_i1 (.D(SLO[0]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i1.GSR = "DISABLED";
    FD1P3AX SLO_i2 (.D(SLO[1]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i2.GSR = "DISABLED";
    FD1P3AX SLO_i3 (.D(SLO[2]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i3.GSR = "DISABLED";
    FD1P3AX SLO_i4 (.D(SLO[3]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i4.GSR = "DISABLED";
    FD1P3AX SLO_i5 (.D(SLO[4]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i5.GSR = "DISABLED";
    FD1P3AX SLO_i6 (.D(SLO[5]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i6.GSR = "DISABLED";
    FD1P3AX SLO_i7 (.D(SLO[6]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i7.GSR = "DISABLED";
    FD1P3AX SLO_i8 (.D(SLO[7]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i8.GSR = "DISABLED";
    FD1P3AX SLO_i9 (.D(SLO[8]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i9.GSR = "DISABLED";
    FD1P3AX SLO_i10 (.D(SLO[9]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i10.GSR = "DISABLED";
    FD1P3AX SLO_i11 (.D(SLO[10]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i11.GSR = "DISABLED";
    FD1P3AX SLO_i12 (.D(SLO[11]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i12.GSR = "DISABLED";
    FD1P3AX SLO_i13 (.D(SLO[12]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i13.GSR = "DISABLED";
    FD1P3AX SLO_i14 (.D(SLO[13]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i14.GSR = "DISABLED";
    FD1P3AX SLO_i15 (.D(SLO[14]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i15.GSR = "DISABLED";
    FD1P3AX SLO_i16 (.D(SLO[15]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i16.GSR = "DISABLED";
    FD1P3AX SLO_i17 (.D(SLO[16]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i17.GSR = "DISABLED";
    FD1P3AX SLO_i18 (.D(SLO[17]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i18.GSR = "DISABLED";
    FD1P3AX SLO_i19 (.D(SLO[18]), .SP(clk_1MHz_derived_322_enable_20), .CK(clk_1MHz_derived_322), 
            .Q(SLO[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i19.GSR = "DISABLED";
    FD1P3IX SLO_i20 (.D(SLO[19]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i20.GSR = "DISABLED";
    FD1P3IX SLO_i21 (.D(SLO[20]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i21.GSR = "DISABLED";
    FD1P3IX SLO_i22 (.D(SLO[21]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i22.GSR = "DISABLED";
    FD1P3IX SLO_i23 (.D(SLO[22]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i23.GSR = "DISABLED";
    FD1P3IX SLO_i24 (.D(SLO[23]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i24.GSR = "DISABLED";
    FD1P3IX SLO_i25 (.D(SLO[24]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i25.GSR = "DISABLED";
    FD1P3IX SLO_i26 (.D(SLO[25]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i26.GSR = "DISABLED";
    FD1P3IX SLO_i27 (.D(SLO[26]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i27.GSR = "DISABLED";
    FD1P3IX SLO_i28 (.D(SLO[27]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i28.GSR = "DISABLED";
    FD1P3IX SLO_i29 (.D(SLO[28]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i29.GSR = "DISABLED";
    FD1P3IX SLO_i30 (.D(SLO[29]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i30.GSR = "DISABLED";
    FD1P3IX SLO_i31 (.D(SLO[30]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i31.GSR = "DISABLED";
    FD1P3IX SLO_i32 (.D(SLO[31]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i32.GSR = "DISABLED";
    FD1P3IX SLO_i33 (.D(SLO[32]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i33.GSR = "DISABLED";
    FD1P3IX SLO_i34 (.D(SLO[33]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i34.GSR = "DISABLED";
    FD1P3IX SLO_i35 (.D(SLO[34]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i35.GSR = "DISABLED";
    FD1P3IX SLO_i36 (.D(SLO[35]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i36.GSR = "DISABLED";
    FD1P3IX SLO_i37 (.D(SLO[36]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i37.GSR = "DISABLED";
    FD1P3IX SLO_i38 (.D(SLO[37]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i38.GSR = "DISABLED";
    FD1P3IX SLO_i39 (.D(SLO[38]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i39.GSR = "DISABLED";
    FD1P3IX SLO_i40 (.D(SLO[39]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i40.GSR = "DISABLED";
    FD1P3IX SLO_i41 (.D(SLO[40]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i41.GSR = "DISABLED";
    FD1P3IX SLO_i42 (.D(SLO[41]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i42.GSR = "DISABLED";
    FD1P3IX SLO_i43 (.D(SLO[42]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i43.GSR = "DISABLED";
    FD1P3IX SLO_i44 (.D(SLO[43]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i44.GSR = "DISABLED";
    FD1P3IX SLO_i45 (.D(SLO[44]), .SP(clk_1MHz_derived_322_enable_46), .CD(MA_Temp_N_5983), 
            .CK(clk_1MHz_derived_322), .Q(SLO[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i45.GSR = "DISABLED";
    LUT4 Select_4070_i21_2_lut (.A(\spi_data_out_r_39__N_5513[16] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6844)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4070_i21_2_lut.init = 16'h8888;
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_6114[1] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_6114[2] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_5852[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_6114[3] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_6114[4] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_6114[5] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_6114[6] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_6114[7] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_6114[8] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_6114[9] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_6114[10] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_6114[11] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_6114[12] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_6114[13] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_6114[14] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_6114[15] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i16 (.D(SLO_buf[30]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i17 (.D(SLO_buf[31]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i18 (.D(SLO_buf[32]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i19 (.D(SLO_buf[33]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i20 (.D(SLO_buf[34]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i21 (.D(SLO_buf[35]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i22 (.D(SLO_buf[36]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i23 (.D(SLO_buf[37]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i24 (.D(SLO_buf[38]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i25 (.D(SLO_buf[39]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i26 (.D(SLO_buf[40]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i27 (.D(SLO_buf[41]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i28 (.D(SLO_buf[42]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i29 (.D(SLO_buf[43]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i30 (.D(SLO_buf[44]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i31 (.D(SLO_buf[45]), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_6114[32] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i33 (.D(\spi_data_out_r_39__N_6114[33] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i33.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i34 (.D(\spi_data_out_r_39__N_6114[34] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i34.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i35 (.D(\spi_data_out_r_39__N_6114[35] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5852[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i35.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i36 (.D(\SLO_buf[10] ), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i36.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i37 (.D(\SLO_buf[11] ), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i37.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i38 (.D(\SLO_buf[12] ), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i38.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i39 (.D(\SLO_buf[13] ), .CK(clk), .CD(n29076), 
            .Q(spi_data_out_r_39__N_5852[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i39.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i1 (.D(n1290[1]), .SP(clk_1MHz_enable_367), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i1.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i2 (.D(n1290[2]), .SP(clk_1MHz_enable_367), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i2.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i3 (.D(n1290[3]), .SP(clk_1MHz_enable_367), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i3.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i4 (.D(n1290[4]), .SP(clk_1MHz_enable_367), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i4.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i5 (.D(n1290[5]), .SP(clk_1MHz_enable_367), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i5.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i6 (.D(n1290[6]), .SP(clk_1MHz_enable_367), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i6.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i7 (.D(n1290[7]), .SP(clk_1MHz_enable_367), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i7.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i8 (.D(n1290[8]), .SP(clk_1MHz_enable_367), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i8.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i9 (.D(n1290[9]), .SP(clk_1MHz_enable_367), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i9.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i10 (.D(n1290[10]), .SP(clk_1MHz_enable_367), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i10.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i11 (.D(n1290[11]), .SP(clk_1MHz_enable_367), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i11.GSR = "DISABLED";
    FD1P3IX Cnt__i1 (.D(n199[1]), .SP(clk_1MHz_enable_374), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i1.GSR = "DISABLED";
    FD1P3IX Cnt__i2 (.D(n199[2]), .SP(clk_1MHz_enable_374), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i3 (.D(n199[3]), .SP(clk_1MHz_enable_374), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i3.GSR = "DISABLED";
    FD1P3IX Cnt__i4 (.D(n199[4]), .SP(clk_1MHz_enable_374), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i4.GSR = "DISABLED";
    FD1P3IX Cnt__i5 (.D(n199[5]), .SP(clk_1MHz_enable_374), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i5.GSR = "DISABLED";
    FD1P3IX Cnt__i6 (.D(n199[6]), .SP(clk_1MHz_enable_374), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i6.GSR = "DISABLED";
    FD1P3IX Cnt__i7 (.D(n199[7]), .SP(clk_1MHz_enable_374), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i7.GSR = "DISABLED";
    LUT4 Select_4070_i18_2_lut (.A(\spi_data_out_r_39__N_4496[16] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6910)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4070_i18_2_lut.init = 16'h8888;
    LUT4 Select_4084_i8_2_lut (.A(\spi_data_out_r_39__N_2338[2] ), .B(spi_data_out_r_39__N_2378), 
         .Z(n8)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4084_i8_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_671 (.A(Cnt_NSL[11]), .B(Cnt_NSL[9]), .C(Cnt_NSL[10]), 
         .D(n4_adj_6918), .Z(n19401)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_671.init = 16'ha080;
    LUT4 Select_4084_i15_2_lut (.A(\spi_data_out_r_39__N_2998[2] ), .B(clear_intrpt_adj_172), 
         .Z(n15)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4084_i15_2_lut.init = 16'h8888;
    LUT4 Select_4084_i11_2_lut (.A(\spi_data_out_r_39__N_2714[2] ), .B(clear_intrpt_adj_173), 
         .Z(n11)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4084_i11_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_672 (.A(Cnt_NSL[7]), .B(Cnt_NSL[8]), .Z(n4_adj_6918)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_672.init = 16'heeee;
    LUT4 Select_4084_i19_2_lut (.A(\spi_data_out_r_39__N_4835[2] ), .B(spi_data_out_r_39__N_4875), 
         .Z(n19)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4084_i19_2_lut.init = 16'h8888;
    CCU2D add_552_7 (.A0(Cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25037), 
          .COUT(n25038), .S0(n153[5]), .S1(n153[6]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_7.INIT0 = 16'h5aaa;
    defparam add_552_7.INIT1 = 16'h5aaa;
    defparam add_552_7.INJECT1_0 = "NO";
    defparam add_552_7.INJECT1_1 = "NO";
    CCU2D add_552_5 (.A0(Cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25036), 
          .COUT(n25037), .S0(n153[3]), .S1(n153[4]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_5.INIT0 = 16'h5aaa;
    defparam add_552_5.INIT1 = 16'h5aaa;
    defparam add_552_5.INJECT1_0 = "NO";
    defparam add_552_5.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_673 (.A(n29275), .B(Cnt[5]), .C(n13378), .D(n19465), 
         .Z(n19439)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i2_4_lut_adj_673.init = 16'hfefa;
    LUT4 i3_4_lut_adj_674 (.A(n19465), .B(Cnt[5]), .C(n29195), .D(n29275), 
         .Z(n19545)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_674.init = 16'hfffe;
    LUT4 i13902_2_lut_3_lut (.A(n19439), .B(n19545), .C(n153[5]), .Z(n199[5])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13902_2_lut_3_lut.init = 16'h7070;
    LUT4 i14525_4_lut (.A(Cnt[0]), .B(Cnt[4]), .C(n27387), .D(Cnt[1]), 
         .Z(n19465)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i14525_4_lut.init = 16'hc8c0;
    LUT4 i10_4_lut_adj_675 (.A(\spi_data_out_r_39__N_3818[16] ), .B(n20_adj_6921), 
         .C(n5_adj_6922), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_6911)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_675.init = 16'hfefc;
    LUT4 Select_4086_i17_2_lut (.A(\spi_data_out_r_39__N_4157[0] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4086_i17_2_lut.init = 16'h8888;
    CCU2D add_552_3 (.A0(Cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25035), 
          .COUT(n25036), .S0(n153[1]), .S1(n153[2]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_3.INIT0 = 16'h5aaa;
    defparam add_552_3.INIT1 = 16'h5aaa;
    defparam add_552_3.INJECT1_0 = "NO";
    defparam add_552_3.INJECT1_1 = "NO";
    LUT4 Select_4086_i3_2_lut (.A(\spi_data_out_r_39__N_1168[0] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4086_i3_2_lut.init = 16'h8888;
    LUT4 Select_4086_i20_2_lut (.A(\spi_data_out_r_39__N_5174[0] ), .B(spi_data_out_r_39__N_5214), 
         .Z(n20)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4086_i20_2_lut.init = 16'h8888;
    LUT4 Select_4086_i15_2_lut (.A(\spi_data_out_r_39__N_2998[0] ), .B(clear_intrpt_adj_172), 
         .Z(n15_adj_174)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4086_i15_2_lut.init = 16'h8888;
    CCU2D add_552_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n25035), 
          .S1(n153[0]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_1.INIT0 = 16'hF000;
    defparam add_552_1.INIT1 = 16'h5555;
    defparam add_552_1.INJECT1_0 = "NO";
    defparam add_552_1.INJECT1_1 = "NO";
    LUT4 Select_4086_i2_2_lut (.A(\spi_data_out_r_39__N_934[0] ), .B(spi_data_out_r_39__N_974), 
         .Z(n2)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4086_i2_2_lut.init = 16'h8888;
    LUT4 Select_4086_i21_2_lut (.A(\spi_data_out_r_39__N_5513[0] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4086_i21_2_lut.init = 16'h8888;
    LUT4 Select_4086_i4_2_lut (.A(\spi_data_out_r_39__N_1402[0] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_175)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4086_i4_2_lut.init = 16'h8888;
    LUT4 Select_4086_i11_2_lut (.A(\spi_data_out_r_39__N_2714[0] ), .B(clear_intrpt_adj_173), 
         .Z(n11_adj_176)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4086_i11_2_lut.init = 16'h8888;
    LUT4 n19439_bdd_3_lut_23072 (.A(n19439), .B(n19545), .C(MA_Temp), 
         .Z(n28794)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam n19439_bdd_3_lut_23072.init = 16'h7070;
    LUT4 i20_4_lut (.A(n27), .B(n40), .C(n36), .D(n28), .Z(\spi_data_out_r[1] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i6_4_lut_adj_676 (.A(\spi_data_out_r_39__N_2643[1] ), .B(\spi_data_out_r_39__N_2856[1] ), 
         .C(clear_intrpt_adj_177), .D(clear_intrpt), .Z(n27)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_676.init = 16'heca0;
    LUT4 i19_4_lut (.A(n31), .B(n38), .C(n4_adj_6931), .D(n22_adj_6932), 
         .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i15_4_lut (.A(\spi_data_out_r_39__N_934[1] ), .B(n30), .C(n19_adj_6933), 
         .D(spi_data_out_r_39__N_974), .Z(n36)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i15_4_lut.init = 16'hfefc;
    LUT4 i7_4_lut (.A(\spi_data_out_r_39__N_4157[1] ), .B(\spi_data_out_r_39__N_1168[1] ), 
         .C(spi_data_out_r_39__N_4197), .D(spi_data_out_r_39__N_1208), .Z(n28)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i7_4_lut.init = 16'heca0;
    LUT4 i10_4_lut_adj_677 (.A(\spi_data_out_r_39__N_2927[1] ), .B(\spi_data_out_r_39__N_2785[1] ), 
         .C(clear_intrpt_adj_178), .D(clear_intrpt_adj_179), .Z(n31)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i10_4_lut_adj_677.init = 16'heca0;
    LUT4 i17_4_lut (.A(n8_adj_6936), .B(n34), .C(n24_adj_6937), .D(n15_adj_6938), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 Select_4085_i4_2_lut (.A(\spi_data_out_r_39__N_1402[1] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6931)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4085_i4_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_678 (.A(\spi_data_out_r_39__N_5174[1] ), .B(\spi_data_out_r_39__N_3818[1] ), 
         .C(spi_data_out_r_39__N_5214), .D(spi_data_out_r_39__N_3858), .Z(n22_adj_6932)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_678.init = 16'heca0;
    LUT4 Select_4085_i8_2_lut (.A(\spi_data_out_r_39__N_2338[1] ), .B(spi_data_out_r_39__N_2378), 
         .Z(n8_adj_6936)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4085_i8_2_lut.init = 16'h8888;
    LUT4 n19439_bdd_4_lut_23207 (.A(n19439), .B(n29271), .C(MA_Temp), 
         .D(Cnt[5]), .Z(n28795)) /* synthesis lut_function=(!(A+!(B (C)+!B !(C (D)+!C !(D))))) */ ;
    defparam n19439_bdd_4_lut_23207.init = 16'h4150;
    LUT4 Select_4065_i18_2_lut (.A(\spi_data_out_r_39__N_4496[21] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6939)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4065_i18_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_679 (.A(spi_data_out_r_39__N_5852[1]), .B(n26_adj_6940), 
         .C(n11_adj_6941), .D(spi_data_out_r_39__N_5892), .Z(n34)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i13_4_lut_adj_679.init = 16'hfefc;
    LUT4 i3_4_lut_adj_680 (.A(\spi_data_out_r_39__N_4496[1] ), .B(\spi_data_out_r_39__N_1870[1] ), 
         .C(spi_data_out_r_39__N_4536), .D(spi_data_out_r_39__N_1910), .Z(n24_adj_6937)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_680.init = 16'heca0;
    LUT4 Select_4085_i15_2_lut (.A(\spi_data_out_r_39__N_2998[1] ), .B(clear_intrpt_adj_172), 
         .Z(n15_adj_6938)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4085_i15_2_lut.init = 16'h8888;
    LUT4 i9_4_lut (.A(\spi_data_out_r_39__N_2104[1] ), .B(\spi_data_out_r_39__N_2572[1] ), 
         .C(spi_data_out_r_39__N_2144), .D(clear_intrpt_adj_180), .Z(n30)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i9_4_lut.init = 16'heca0;
    LUT4 Select_4085_i19_2_lut (.A(\spi_data_out_r_39__N_4835[1] ), .B(spi_data_out_r_39__N_4875), 
         .Z(n19_adj_6933)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4085_i19_2_lut.init = 16'h8888;
    LUT4 i5_4_lut_adj_681 (.A(\spi_data_out_r_39__N_5513[1] ), .B(\spi_data_out_r_39__N_1636[1] ), 
         .C(spi_data_out_r_39__N_5553), .D(spi_data_out_r_39__N_1676), .Z(n26_adj_6940)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i5_4_lut_adj_681.init = 16'heca0;
    LUT4 Select_4085_i11_2_lut (.A(\spi_data_out_r_39__N_2714[1] ), .B(clear_intrpt_adj_173), 
         .Z(n11_adj_6941)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4085_i11_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_682 (.A(n3_adj_6943), .B(n26_adj_6944), .C(n22_adj_6945), 
         .D(n21_adj_6946), .Z(\spi_data_out_r[3] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_682.init = 16'hfffe;
    LUT4 Select_4083_i3_2_lut (.A(\spi_data_out_r_39__N_1168[3] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_6943)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4083_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_683 (.A(n18_adj_6947), .B(n24_adj_6948), .C(n18_adj_6949), 
         .D(n4_adj_6950), .Z(n26_adj_6944)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_683.init = 16'hfffe;
    LUT4 i8_4_lut_adj_684 (.A(\spi_data_out_r_39__N_4835[3] ), .B(n16_adj_6951), 
         .C(n17_adj_6952), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6945)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_684.init = 16'hfefc;
    LUT4 Select_4083_i21_2_lut (.A(\spi_data_out_r_39__N_5513[3] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6946)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4083_i21_2_lut.init = 16'h8888;
    LUT4 n28797_bdd_3_lut (.A(n28797), .B(n28794), .C(n29192), .Z(MA_Temp_N_5972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28797_bdd_3_lut.init = 16'hcaca;
    LUT4 Select_4083_i18_2_lut (.A(\spi_data_out_r_39__N_4496[3] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6947)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4083_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_685 (.A(\spi_data_out_r_39__N_3818[3] ), .B(n20_adj_6953), 
         .C(n5_adj_6954), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_6948)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_685.init = 16'hfefc;
    LUT4 i4_4_lut_adj_686 (.A(\spi_data_out_r_39__N_2104[3] ), .B(\spi_data_out_r_39__N_1870[3] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6949)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_686.init = 16'heca0;
    LUT4 Select_4083_i4_2_lut (.A(\spi_data_out_r_39__N_1402[3] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6950)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4083_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_687 (.A(\spi_data_out_r_39__N_2338[3] ), .B(\spi_data_out_r_39__N_5174[3] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_6953)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_687.init = 16'heca0;
    LUT4 Select_4083_i5_2_lut (.A(\spi_data_out_r_39__N_1636[3] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6954)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4083_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_688 (.A(\spi_data_out_r_39__N_934[3] ), .B(spi_data_out_r_39__N_5852[3]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6951)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_688.init = 16'heca0;
    LUT4 Select_4083_i17_2_lut (.A(\spi_data_out_r_39__N_4157[3] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6952)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4083_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_689 (.A(n3_adj_6955), .B(n26_adj_6956), .C(n22_adj_6957), 
         .D(n21_adj_6958), .Z(\spi_data_out_r[4] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_689.init = 16'hfffe;
    LUT4 Select_4082_i3_2_lut (.A(\spi_data_out_r_39__N_1168[4] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_6955)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4082_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_690 (.A(n18_adj_6959), .B(n24_adj_6960), .C(n18_adj_6961), 
         .D(n4_adj_6962), .Z(n26_adj_6956)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_690.init = 16'hfffe;
    LUT4 i8_4_lut_adj_691 (.A(\spi_data_out_r_39__N_4835[4] ), .B(n16_adj_6963), 
         .C(n17_adj_6964), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6957)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_691.init = 16'hfefc;
    LUT4 Select_4082_i21_2_lut (.A(\spi_data_out_r_39__N_5513[4] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6958)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4082_i21_2_lut.init = 16'h8888;
    LUT4 Select_4082_i18_2_lut (.A(\spi_data_out_r_39__N_4496[4] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6959)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4082_i18_2_lut.init = 16'h8888;
    LUT4 i4_4_lut_adj_692 (.A(\spi_data_out_r_39__N_2104[16] ), .B(\spi_data_out_r_39__N_1870[16] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6912)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_692.init = 16'heca0;
    LUT4 i10_4_lut_adj_693 (.A(\spi_data_out_r_39__N_3818[4] ), .B(n20_adj_6965), 
         .C(n5_adj_6966), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_6960)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_693.init = 16'hfefc;
    LUT4 i4_4_lut_adj_694 (.A(\spi_data_out_r_39__N_2104[4] ), .B(\spi_data_out_r_39__N_1870[4] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6961)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_694.init = 16'heca0;
    LUT4 Select_4070_i4_2_lut (.A(\spi_data_out_r_39__N_1402[16] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6913)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4070_i4_2_lut.init = 16'h8888;
    LUT4 Select_4082_i4_2_lut (.A(\spi_data_out_r_39__N_1402[4] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6962)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4082_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_695 (.A(\spi_data_out_r_39__N_2338[4] ), .B(\spi_data_out_r_39__N_5174[4] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_6965)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_695.init = 16'heca0;
    LUT4 Select_4082_i5_2_lut (.A(\spi_data_out_r_39__N_1636[4] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6966)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4082_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_696 (.A(\spi_data_out_r_39__N_934[4] ), .B(spi_data_out_r_39__N_5852[4]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6963)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_696.init = 16'heca0;
    LUT4 Select_4082_i17_2_lut (.A(\spi_data_out_r_39__N_4157[4] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6964)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4082_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_697 (.A(n3_adj_6967), .B(n26_adj_6968), .C(n22_adj_6969), 
         .D(n21_adj_6970), .Z(\spi_data_out_r[5] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_697.init = 16'hfffe;
    LUT4 Select_4081_i3_2_lut (.A(\spi_data_out_r_39__N_1168[5] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_6967)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4081_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_698 (.A(n18_adj_6971), .B(n24_adj_6972), .C(n18_adj_6973), 
         .D(n4_adj_6974), .Z(n26_adj_6968)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_698.init = 16'hfffe;
    LUT4 i8_4_lut_adj_699 (.A(\spi_data_out_r_39__N_4835[5] ), .B(n16_adj_6975), 
         .C(n17_adj_6976), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6969)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_699.init = 16'hfefc;
    LUT4 Select_4081_i21_2_lut (.A(\spi_data_out_r_39__N_5513[5] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6970)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4081_i21_2_lut.init = 16'h8888;
    LUT4 Select_4081_i18_2_lut (.A(\spi_data_out_r_39__N_4496[5] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6971)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4081_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_700 (.A(\spi_data_out_r_39__N_3818[5] ), .B(n20_adj_6977), 
         .C(n5_adj_6978), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_6972)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_700.init = 16'hfefc;
    LUT4 i4_4_lut_adj_701 (.A(\spi_data_out_r_39__N_2104[5] ), .B(\spi_data_out_r_39__N_1870[5] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6973)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_701.init = 16'heca0;
    LUT4 Select_4081_i4_2_lut (.A(\spi_data_out_r_39__N_1402[5] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6974)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4081_i4_2_lut.init = 16'h8888;
    FD1P3IX MA_Temp_474 (.D(MA_Temp_N_5972), .SP(clk_1MHz_enable_377), .CD(n29239), 
            .CK(clk_1MHz), .Q(MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam MA_Temp_474.GSR = "DISABLED";
    LUT4 i6_4_lut_adj_702 (.A(\spi_data_out_r_39__N_2338[5] ), .B(\spi_data_out_r_39__N_5174[5] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_6977)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_702.init = 16'heca0;
    LUT4 Select_4081_i5_2_lut (.A(\spi_data_out_r_39__N_1636[5] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6978)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4081_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_703 (.A(\spi_data_out_r_39__N_934[5] ), .B(spi_data_out_r_39__N_5852[5]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6975)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_703.init = 16'heca0;
    LUT4 Select_4081_i17_2_lut (.A(\spi_data_out_r_39__N_4157[5] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6976)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4081_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_704 (.A(n3_adj_6979), .B(n26_adj_6980), .C(n22_adj_6981), 
         .D(n21_adj_6982), .Z(\spi_data_out_r[6] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_704.init = 16'hfffe;
    LUT4 Select_4080_i3_2_lut (.A(\spi_data_out_r_39__N_1168[6] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_6979)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4080_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_705 (.A(n18_adj_6983), .B(n24_adj_6984), .C(n18_adj_6985), 
         .D(n4_adj_6986), .Z(n26_adj_6980)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_705.init = 16'hfffe;
    LUT4 i8_4_lut_adj_706 (.A(\spi_data_out_r_39__N_4835[6] ), .B(n16_adj_6987), 
         .C(n17_adj_6988), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6981)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_706.init = 16'hfefc;
    LUT4 Select_4080_i21_2_lut (.A(\spi_data_out_r_39__N_5513[6] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6982)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4080_i21_2_lut.init = 16'h8888;
    LUT4 Select_4080_i18_2_lut (.A(\spi_data_out_r_39__N_4496[6] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6983)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4080_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_707 (.A(\spi_data_out_r_39__N_3818[6] ), .B(n20_adj_6989), 
         .C(n5_adj_6990), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_6984)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_707.init = 16'hfefc;
    LUT4 i4_4_lut_adj_708 (.A(\spi_data_out_r_39__N_2104[6] ), .B(\spi_data_out_r_39__N_1870[6] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6985)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_708.init = 16'heca0;
    LUT4 Select_4080_i4_2_lut (.A(\spi_data_out_r_39__N_1402[6] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6986)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4080_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_709 (.A(\spi_data_out_r_39__N_2338[6] ), .B(\spi_data_out_r_39__N_5174[6] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_6989)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_709.init = 16'heca0;
    LUT4 Select_4080_i5_2_lut (.A(\spi_data_out_r_39__N_1636[6] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6990)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4080_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_710 (.A(\spi_data_out_r_39__N_934[6] ), .B(spi_data_out_r_39__N_5852[6]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6987)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_710.init = 16'heca0;
    LUT4 Select_4080_i17_2_lut (.A(\spi_data_out_r_39__N_4157[6] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6988)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4080_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_711 (.A(n3_adj_6991), .B(n26_adj_6992), .C(n22_adj_6993), 
         .D(n21_adj_6994), .Z(\spi_data_out_r[7] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_711.init = 16'hfffe;
    LUT4 Select_4079_i3_2_lut (.A(\spi_data_out_r_39__N_1168[7] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_6991)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4079_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_712 (.A(n18_adj_6995), .B(n24_adj_6996), .C(n18_adj_6997), 
         .D(n4_adj_6998), .Z(n26_adj_6992)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_712.init = 16'hfffe;
    LUT4 i8_4_lut_adj_713 (.A(\spi_data_out_r_39__N_4835[7] ), .B(n16_adj_6999), 
         .C(n17_adj_7000), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_6993)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_713.init = 16'hfefc;
    LUT4 Select_4079_i21_2_lut (.A(\spi_data_out_r_39__N_5513[7] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_6994)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4079_i21_2_lut.init = 16'h8888;
    LUT4 Select_4079_i18_2_lut (.A(\spi_data_out_r_39__N_4496[7] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_6995)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4079_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_714 (.A(\spi_data_out_r_39__N_3818[7] ), .B(n20_adj_7001), 
         .C(n5_adj_7002), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_6996)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_714.init = 16'hfefc;
    LUT4 i4_4_lut_adj_715 (.A(\spi_data_out_r_39__N_2104[7] ), .B(\spi_data_out_r_39__N_1870[7] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_6997)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_715.init = 16'heca0;
    LUT4 Select_4079_i4_2_lut (.A(\spi_data_out_r_39__N_1402[7] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_6998)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4079_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_716 (.A(\spi_data_out_r_39__N_2338[7] ), .B(\spi_data_out_r_39__N_5174[7] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_7001)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_716.init = 16'heca0;
    LUT4 Select_4079_i5_2_lut (.A(\spi_data_out_r_39__N_1636[7] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_7002)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4079_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_717 (.A(\spi_data_out_r_39__N_934[7] ), .B(spi_data_out_r_39__N_5852[7]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6999)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_717.init = 16'heca0;
    LUT4 Select_4079_i17_2_lut (.A(\spi_data_out_r_39__N_4157[7] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_7000)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4079_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_718 (.A(n3_adj_7003), .B(n26_adj_7004), .C(n22_adj_7005), 
         .D(n21_adj_7006), .Z(\spi_data_out_r[8] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_718.init = 16'hfffe;
    LUT4 Select_4078_i3_2_lut (.A(\spi_data_out_r_39__N_1168[8] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_7003)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4078_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_719 (.A(n18_adj_7007), .B(n24_adj_7008), .C(n18_adj_7009), 
         .D(n4_adj_7010), .Z(n26_adj_7004)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_719.init = 16'hfffe;
    LUT4 i8_4_lut_adj_720 (.A(\spi_data_out_r_39__N_4835[8] ), .B(n16_adj_7011), 
         .C(n17_adj_7012), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_7005)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_720.init = 16'hfefc;
    LUT4 Select_4078_i21_2_lut (.A(\spi_data_out_r_39__N_5513[8] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_7006)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4078_i21_2_lut.init = 16'h8888;
    LUT4 Select_4078_i18_2_lut (.A(\spi_data_out_r_39__N_4496[8] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_7007)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4078_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_721 (.A(\spi_data_out_r_39__N_3818[8] ), .B(n20_adj_7013), 
         .C(n5_adj_7014), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_7008)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_721.init = 16'hfefc;
    LUT4 i4_4_lut_adj_722 (.A(\spi_data_out_r_39__N_2104[8] ), .B(\spi_data_out_r_39__N_1870[8] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_7009)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_722.init = 16'heca0;
    LUT4 Select_4078_i4_2_lut (.A(\spi_data_out_r_39__N_1402[8] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_7010)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4078_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_723 (.A(\spi_data_out_r_39__N_2338[8] ), .B(\spi_data_out_r_39__N_5174[8] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_7013)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_723.init = 16'heca0;
    LUT4 Select_4078_i5_2_lut (.A(\spi_data_out_r_39__N_1636[8] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_7014)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4078_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_724 (.A(\spi_data_out_r_39__N_934[8] ), .B(spi_data_out_r_39__N_5852[8]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_7011)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_724.init = 16'heca0;
    LUT4 Select_4078_i17_2_lut (.A(\spi_data_out_r_39__N_4157[8] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_7012)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4078_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_725 (.A(n3_adj_7015), .B(n26_adj_7016), .C(n22_adj_7017), 
         .D(n21_adj_7018), .Z(\spi_data_out_r[9] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_725.init = 16'hfffe;
    LUT4 Select_4077_i3_2_lut (.A(\spi_data_out_r_39__N_1168[9] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_7015)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4077_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_726 (.A(n18_adj_7019), .B(n24_adj_7020), .C(n18_adj_7021), 
         .D(n4_adj_7022), .Z(n26_adj_7016)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_726.init = 16'hfffe;
    LUT4 i8_4_lut_adj_727 (.A(\spi_data_out_r_39__N_4835[9] ), .B(n16_adj_7023), 
         .C(n17_adj_7024), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_7017)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_727.init = 16'hfefc;
    LUT4 Select_4077_i21_2_lut (.A(\spi_data_out_r_39__N_5513[9] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_7018)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4077_i21_2_lut.init = 16'h8888;
    LUT4 Select_4077_i18_2_lut (.A(\spi_data_out_r_39__N_4496[9] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_7019)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4077_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_728 (.A(\spi_data_out_r_39__N_3818[9] ), .B(n20_adj_7025), 
         .C(n5_adj_7026), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_7020)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_728.init = 16'hfefc;
    LUT4 i4_4_lut_adj_729 (.A(\spi_data_out_r_39__N_2104[9] ), .B(\spi_data_out_r_39__N_1870[9] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_7021)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_729.init = 16'heca0;
    LUT4 Select_4077_i4_2_lut (.A(\spi_data_out_r_39__N_1402[9] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_7022)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4077_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_730 (.A(\spi_data_out_r_39__N_2338[9] ), .B(\spi_data_out_r_39__N_5174[9] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_7025)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_730.init = 16'heca0;
    LUT4 Select_4077_i5_2_lut (.A(\spi_data_out_r_39__N_1636[9] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_7026)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4077_i5_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_731 (.A(\spi_data_out_r_39__N_2338[16] ), .B(\spi_data_out_r_39__N_5174[16] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_6921)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_731.init = 16'heca0;
    LUT4 i2_4_lut_adj_732 (.A(\spi_data_out_r_39__N_934[9] ), .B(spi_data_out_r_39__N_5852[9]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_7023)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_732.init = 16'heca0;
    LUT4 Select_4077_i17_2_lut (.A(\spi_data_out_r_39__N_4157[9] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_7024)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4077_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_733 (.A(n3_adj_7027), .B(n26_adj_7028), .C(n22_adj_7029), 
         .D(n21_adj_7030), .Z(\spi_data_out_r[10] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_733.init = 16'hfffe;
    LUT4 Select_4076_i3_2_lut (.A(\spi_data_out_r_39__N_1168[10] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_7027)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4076_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_734 (.A(n18_adj_7031), .B(n24_adj_7032), .C(n18_adj_7033), 
         .D(n4_adj_7034), .Z(n26_adj_7028)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_734.init = 16'hfffe;
    LUT4 i8_4_lut_adj_735 (.A(\spi_data_out_r_39__N_4835[10] ), .B(n16_adj_7035), 
         .C(n17_adj_7036), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_7029)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_735.init = 16'hfefc;
    LUT4 Select_4076_i21_2_lut (.A(\spi_data_out_r_39__N_5513[10] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_7030)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4076_i21_2_lut.init = 16'h8888;
    LUT4 Select_4076_i18_2_lut (.A(\spi_data_out_r_39__N_4496[10] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_7031)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4076_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_736 (.A(\spi_data_out_r_39__N_3818[10] ), .B(n20_adj_7037), 
         .C(n5_adj_7038), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_7032)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_736.init = 16'hfefc;
    LUT4 i4_4_lut_adj_737 (.A(\spi_data_out_r_39__N_2104[10] ), .B(\spi_data_out_r_39__N_1870[10] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_7033)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_737.init = 16'heca0;
    LUT4 Select_4076_i4_2_lut (.A(\spi_data_out_r_39__N_1402[10] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_7034)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4076_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_738 (.A(\spi_data_out_r_39__N_2338[10] ), .B(\spi_data_out_r_39__N_5174[10] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_7037)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_738.init = 16'heca0;
    LUT4 Select_4076_i5_2_lut (.A(\spi_data_out_r_39__N_1636[10] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_7038)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4076_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_739 (.A(\spi_data_out_r_39__N_934[10] ), .B(spi_data_out_r_39__N_5852[10]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_7035)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_739.init = 16'heca0;
    LUT4 Select_4076_i17_2_lut (.A(\spi_data_out_r_39__N_4157[10] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_7036)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4076_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_740 (.A(n3_adj_7039), .B(n26_adj_7040), .C(n22_adj_7041), 
         .D(n21_adj_7042), .Z(\spi_data_out_r[11] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_740.init = 16'hfffe;
    LUT4 Select_4075_i3_2_lut (.A(\spi_data_out_r_39__N_1168[11] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_7039)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4075_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_741 (.A(n18_adj_7043), .B(n24_adj_7044), .C(n18_adj_7045), 
         .D(n4_adj_7046), .Z(n26_adj_7040)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_741.init = 16'hfffe;
    LUT4 i8_4_lut_adj_742 (.A(\spi_data_out_r_39__N_4835[11] ), .B(n16_adj_7047), 
         .C(n17_adj_7048), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_7041)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_742.init = 16'hfefc;
    LUT4 Select_4075_i21_2_lut (.A(\spi_data_out_r_39__N_5513[11] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_7042)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4075_i21_2_lut.init = 16'h8888;
    LUT4 Select_4075_i18_2_lut (.A(\spi_data_out_r_39__N_4496[11] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_7043)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4075_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_743 (.A(\spi_data_out_r_39__N_3818[11] ), .B(n20_adj_7049), 
         .C(n5_adj_7050), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_7044)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_743.init = 16'hfefc;
    LUT4 i4_4_lut_adj_744 (.A(\spi_data_out_r_39__N_2104[11] ), .B(\spi_data_out_r_39__N_1870[11] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_7045)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_744.init = 16'heca0;
    LUT4 Select_4075_i4_2_lut (.A(\spi_data_out_r_39__N_1402[11] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_7046)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4075_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_745 (.A(\spi_data_out_r_39__N_2338[11] ), .B(\spi_data_out_r_39__N_5174[11] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_7049)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_745.init = 16'heca0;
    LUT4 Select_4075_i5_2_lut (.A(\spi_data_out_r_39__N_1636[11] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_7050)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4075_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_746 (.A(\spi_data_out_r_39__N_934[11] ), .B(spi_data_out_r_39__N_5852[11]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_7047)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_746.init = 16'heca0;
    LUT4 Select_4075_i17_2_lut (.A(\spi_data_out_r_39__N_4157[11] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_7048)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4075_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_747 (.A(n3_adj_7051), .B(n26_adj_7052), .C(n22_adj_7053), 
         .D(n21_adj_7054), .Z(\spi_data_out_r[12] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_747.init = 16'hfffe;
    LUT4 Select_4074_i3_2_lut (.A(\spi_data_out_r_39__N_1168[12] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_7051)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4074_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_748 (.A(n18_adj_7055), .B(n24_adj_7056), .C(n18_adj_7057), 
         .D(n4_adj_7058), .Z(n26_adj_7052)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_748.init = 16'hfffe;
    LUT4 i8_4_lut_adj_749 (.A(\spi_data_out_r_39__N_4835[12] ), .B(n16_adj_7059), 
         .C(n17_adj_7060), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_7053)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_749.init = 16'hfefc;
    LUT4 Select_4074_i21_2_lut (.A(\spi_data_out_r_39__N_5513[12] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_7054)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4074_i21_2_lut.init = 16'h8888;
    LUT4 Select_4074_i18_2_lut (.A(\spi_data_out_r_39__N_4496[12] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_7055)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4074_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_750 (.A(\spi_data_out_r_39__N_3818[12] ), .B(n20_adj_7061), 
         .C(n5_adj_7062), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_7056)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_750.init = 16'hfefc;
    LUT4 i4_4_lut_adj_751 (.A(\spi_data_out_r_39__N_2104[12] ), .B(\spi_data_out_r_39__N_1870[12] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_7057)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_751.init = 16'heca0;
    LUT4 Select_4074_i4_2_lut (.A(\spi_data_out_r_39__N_1402[12] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_7058)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4074_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_752 (.A(\spi_data_out_r_39__N_2338[12] ), .B(\spi_data_out_r_39__N_5174[12] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_7061)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_752.init = 16'heca0;
    LUT4 Select_4074_i5_2_lut (.A(\spi_data_out_r_39__N_1636[12] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_7062)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4074_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_753 (.A(\spi_data_out_r_39__N_934[12] ), .B(spi_data_out_r_39__N_5852[12]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_7059)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_753.init = 16'heca0;
    LUT4 Select_4074_i17_2_lut (.A(\spi_data_out_r_39__N_4157[12] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_7060)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4074_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_754 (.A(n3_adj_7063), .B(n26_adj_7064), .C(n22_adj_7065), 
         .D(n21_adj_7066), .Z(\spi_data_out_r[13] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_754.init = 16'hfffe;
    LUT4 Select_4073_i3_2_lut (.A(\spi_data_out_r_39__N_1168[13] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_7063)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4073_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_755 (.A(n18_adj_7067), .B(n24_adj_7068), .C(n18_adj_7069), 
         .D(n4_adj_7070), .Z(n26_adj_7064)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_755.init = 16'hfffe;
    LUT4 i8_4_lut_adj_756 (.A(\spi_data_out_r_39__N_4835[13] ), .B(n16_adj_7071), 
         .C(n17_adj_7072), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_7065)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_756.init = 16'hfefc;
    LUT4 Select_4073_i21_2_lut (.A(\spi_data_out_r_39__N_5513[13] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_7066)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4073_i21_2_lut.init = 16'h8888;
    LUT4 Select_4073_i18_2_lut (.A(\spi_data_out_r_39__N_4496[13] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_7067)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4073_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_757 (.A(\spi_data_out_r_39__N_3818[13] ), .B(n20_adj_7073), 
         .C(n5_adj_7074), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_7068)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_757.init = 16'hfefc;
    LUT4 i4_4_lut_adj_758 (.A(\spi_data_out_r_39__N_2104[13] ), .B(\spi_data_out_r_39__N_1870[13] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_7069)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_758.init = 16'heca0;
    LUT4 Select_4073_i4_2_lut (.A(\spi_data_out_r_39__N_1402[13] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_7070)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4073_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_759 (.A(\spi_data_out_r_39__N_2338[13] ), .B(\spi_data_out_r_39__N_5174[13] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_7073)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_759.init = 16'heca0;
    LUT4 Select_4073_i5_2_lut (.A(\spi_data_out_r_39__N_1636[13] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_7074)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4073_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_760 (.A(\spi_data_out_r_39__N_934[13] ), .B(spi_data_out_r_39__N_5852[13]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_7071)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_760.init = 16'heca0;
    LUT4 Select_4073_i17_2_lut (.A(\spi_data_out_r_39__N_4157[13] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_7072)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4073_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_761 (.A(n3_adj_7075), .B(n26_adj_7076), .C(n22_adj_7077), 
         .D(n21_adj_7078), .Z(\spi_data_out_r[14] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_761.init = 16'hfffe;
    LUT4 Select_4072_i3_2_lut (.A(\spi_data_out_r_39__N_1168[14] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_7075)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4072_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_762 (.A(n18_adj_7079), .B(n24_adj_7080), .C(n18_adj_7081), 
         .D(n4_adj_7082), .Z(n26_adj_7076)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_762.init = 16'hfffe;
    LUT4 i8_4_lut_adj_763 (.A(\spi_data_out_r_39__N_4835[14] ), .B(n16_adj_7083), 
         .C(n17_adj_7084), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_7077)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_763.init = 16'hfefc;
    LUT4 Select_4072_i21_2_lut (.A(\spi_data_out_r_39__N_5513[14] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_7078)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4072_i21_2_lut.init = 16'h8888;
    LUT4 Select_4072_i18_2_lut (.A(\spi_data_out_r_39__N_4496[14] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_7079)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4072_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_764 (.A(\spi_data_out_r_39__N_3818[14] ), .B(n20_adj_7085), 
         .C(n5_adj_7086), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_7080)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_764.init = 16'hfefc;
    LUT4 i4_4_lut_adj_765 (.A(\spi_data_out_r_39__N_2104[14] ), .B(\spi_data_out_r_39__N_1870[14] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_7081)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_765.init = 16'heca0;
    LUT4 Select_4072_i4_2_lut (.A(\spi_data_out_r_39__N_1402[14] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_7082)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4072_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_766 (.A(\spi_data_out_r_39__N_2338[14] ), .B(\spi_data_out_r_39__N_5174[14] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_7085)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_766.init = 16'heca0;
    LUT4 Select_4072_i5_2_lut (.A(\spi_data_out_r_39__N_1636[14] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_7086)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4072_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_767 (.A(\spi_data_out_r_39__N_934[14] ), .B(spi_data_out_r_39__N_5852[14]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_7083)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_767.init = 16'heca0;
    LUT4 Select_4072_i17_2_lut (.A(\spi_data_out_r_39__N_4157[14] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_7084)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4072_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_768 (.A(n3_adj_7087), .B(n26_adj_7088), .C(n22_adj_7089), 
         .D(n21_adj_7090), .Z(\spi_data_out_r[15] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_768.init = 16'hfffe;
    LUT4 Select_4071_i3_2_lut (.A(\spi_data_out_r_39__N_1168[15] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_7087)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4071_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_769 (.A(n18_adj_7091), .B(n24_adj_7092), .C(n18_adj_7093), 
         .D(n4_adj_7094), .Z(n26_adj_7088)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_769.init = 16'hfffe;
    LUT4 i8_4_lut_adj_770 (.A(\spi_data_out_r_39__N_4835[15] ), .B(n16_adj_6786), 
         .C(n17_adj_6787), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_7089)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_770.init = 16'hfefc;
    LUT4 Select_4070_i5_2_lut (.A(\spi_data_out_r_39__N_1636[16] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_6922)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4070_i5_2_lut.init = 16'h8888;
    LUT4 Select_4071_i21_2_lut (.A(\spi_data_out_r_39__N_5513[15] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_7090)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4071_i21_2_lut.init = 16'h8888;
    LUT4 Select_4071_i18_2_lut (.A(\spi_data_out_r_39__N_4496[15] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_7091)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4071_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_771 (.A(\spi_data_out_r_39__N_3818[15] ), .B(n20_adj_7095), 
         .C(n5), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_7092)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_771.init = 16'hfefc;
    LUT4 i4_4_lut_adj_772 (.A(\spi_data_out_r_39__N_2104[15] ), .B(\spi_data_out_r_39__N_1870[15] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_7093)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_772.init = 16'heca0;
    LUT4 Select_4071_i4_2_lut (.A(\spi_data_out_r_39__N_1402[15] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_7094)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4071_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_773 (.A(\spi_data_out_r_39__N_2338[15] ), .B(\spi_data_out_r_39__N_5174[15] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_7095)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_773.init = 16'heca0;
    LUT4 i2_4_lut_adj_774 (.A(\spi_data_out_r_39__N_934[16] ), .B(spi_data_out_r_39__N_5852[16]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_6914)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_774.init = 16'heca0;
    LUT4 Select_4070_i17_2_lut (.A(\spi_data_out_r_39__N_4157[16] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_6915)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4070_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_775 (.A(n3_adj_7096), .B(n26_adj_7097), .C(n22_adj_7098), 
         .D(n21_adj_7099), .Z(\spi_data_out_r[17] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_775.init = 16'hfffe;
    LUT4 Select_4069_i3_2_lut (.A(\spi_data_out_r_39__N_1168[17] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_7096)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4069_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_776 (.A(n18_adj_7100), .B(n24_adj_7101), .C(n18_adj_7102), 
         .D(n4_adj_7103), .Z(n26_adj_7097)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_776.init = 16'hfffe;
    LUT4 i8_4_lut_adj_777 (.A(\spi_data_out_r_39__N_4835[17] ), .B(n16_adj_7104), 
         .C(n17_adj_7105), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_7098)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_777.init = 16'hfefc;
    LUT4 Select_4069_i21_2_lut (.A(\spi_data_out_r_39__N_5513[17] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_7099)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4069_i21_2_lut.init = 16'h8888;
    LUT4 Select_4069_i18_2_lut (.A(\spi_data_out_r_39__N_4496[17] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_7100)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4069_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_778 (.A(\spi_data_out_r_39__N_3818[17] ), .B(n20_adj_7106), 
         .C(n5_adj_7107), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_7101)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_778.init = 16'hfefc;
    LUT4 i4_4_lut_adj_779 (.A(\spi_data_out_r_39__N_2104[17] ), .B(\spi_data_out_r_39__N_1870[17] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_7102)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_779.init = 16'heca0;
    LUT4 Select_4069_i4_2_lut (.A(\spi_data_out_r_39__N_1402[17] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_7103)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4069_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_780 (.A(\spi_data_out_r_39__N_2338[17] ), .B(\spi_data_out_r_39__N_5174[17] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_7106)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_780.init = 16'heca0;
    LUT4 Select_4069_i5_2_lut (.A(\spi_data_out_r_39__N_1636[17] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_7107)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4069_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_781 (.A(\spi_data_out_r_39__N_934[17] ), .B(spi_data_out_r_39__N_5852[17]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_7104)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_781.init = 16'heca0;
    LUT4 Select_4069_i17_2_lut (.A(\spi_data_out_r_39__N_4157[17] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_7105)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4069_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_782 (.A(n3_adj_7108), .B(n26_adj_7109), .C(n22_adj_7110), 
         .D(n21_adj_7111), .Z(\spi_data_out_r[18] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_782.init = 16'hfffe;
    LUT4 Select_4068_i3_2_lut (.A(\spi_data_out_r_39__N_1168[18] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_7108)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4068_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_783 (.A(n18_adj_7112), .B(n24_adj_7113), .C(n18_adj_7114), 
         .D(n4_adj_7115), .Z(n26_adj_7109)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_783.init = 16'hfffe;
    LUT4 i8_4_lut_adj_784 (.A(\spi_data_out_r_39__N_4835[18] ), .B(n16_adj_7116), 
         .C(n17_adj_7117), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_7110)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_784.init = 16'hfefc;
    LUT4 Select_4068_i21_2_lut (.A(\spi_data_out_r_39__N_5513[18] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_7111)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4068_i21_2_lut.init = 16'h8888;
    LUT4 Select_4068_i18_2_lut (.A(\spi_data_out_r_39__N_4496[18] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_7112)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4068_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_785 (.A(\spi_data_out_r_39__N_3818[18] ), .B(n20_adj_7118), 
         .C(n5_adj_7119), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_7113)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_785.init = 16'hfefc;
    LUT4 i4_4_lut_adj_786 (.A(\spi_data_out_r_39__N_2104[18] ), .B(\spi_data_out_r_39__N_1870[18] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_7114)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_786.init = 16'heca0;
    LUT4 Select_4068_i4_2_lut (.A(\spi_data_out_r_39__N_1402[18] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_7115)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4068_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_787 (.A(\spi_data_out_r_39__N_2338[18] ), .B(\spi_data_out_r_39__N_5174[18] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_7118)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_787.init = 16'heca0;
    LUT4 Select_4068_i5_2_lut (.A(\spi_data_out_r_39__N_1636[18] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_7119)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4068_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_788 (.A(\spi_data_out_r_39__N_934[18] ), .B(spi_data_out_r_39__N_5852[18]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_7116)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_788.init = 16'heca0;
    LUT4 Select_4068_i17_2_lut (.A(\spi_data_out_r_39__N_4157[18] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_7117)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4068_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_789 (.A(n3_adj_7120), .B(n26_adj_7121), .C(n22_adj_7122), 
         .D(n21_adj_7123), .Z(\spi_data_out_r[19] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_789.init = 16'hfffe;
    LUT4 Select_4067_i3_2_lut (.A(\spi_data_out_r_39__N_1168[19] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_7120)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4067_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_790 (.A(n18_adj_7124), .B(n24_adj_7125), .C(n18_adj_7126), 
         .D(n4_adj_7127), .Z(n26_adj_7121)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_790.init = 16'hfffe;
    LUT4 i8_4_lut_adj_791 (.A(\spi_data_out_r_39__N_4835[19] ), .B(n16_adj_7128), 
         .C(n17_adj_7129), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_7122)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_791.init = 16'hfefc;
    LUT4 Select_4067_i21_2_lut (.A(\spi_data_out_r_39__N_5513[19] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_7123)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4067_i21_2_lut.init = 16'h8888;
    LUT4 Select_4067_i18_2_lut (.A(\spi_data_out_r_39__N_4496[19] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_7124)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4067_i18_2_lut.init = 16'h8888;
    LUT4 i10_4_lut_adj_792 (.A(\spi_data_out_r_39__N_3818[19] ), .B(n20_adj_7130), 
         .C(n5_adj_7131), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_7125)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_792.init = 16'hfefc;
    LUT4 i4_4_lut_adj_793 (.A(\spi_data_out_r_39__N_2104[19] ), .B(\spi_data_out_r_39__N_1870[19] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_7126)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_793.init = 16'heca0;
    LUT4 Select_4067_i4_2_lut (.A(\spi_data_out_r_39__N_1402[19] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_7127)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4067_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_794 (.A(\spi_data_out_r_39__N_2338[19] ), .B(\spi_data_out_r_39__N_5174[19] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_7130)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_794.init = 16'heca0;
    LUT4 Select_4067_i5_2_lut (.A(\spi_data_out_r_39__N_1636[19] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_7131)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4067_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_795 (.A(\spi_data_out_r_39__N_934[19] ), .B(spi_data_out_r_39__N_5852[19]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_7128)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_795.init = 16'heca0;
    LUT4 Select_4067_i17_2_lut (.A(\spi_data_out_r_39__N_4157[19] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_7129)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4067_i17_2_lut.init = 16'h8888;
    LUT4 i13_4_lut_adj_796 (.A(n3_adj_7132), .B(n26_adj_7133), .C(n22_adj_7134), 
         .D(n21_adj_7135), .Z(\spi_data_out_r[20] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_796.init = 16'hfffe;
    LUT4 Select_4066_i3_2_lut (.A(\spi_data_out_r_39__N_1168[20] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_7132)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4066_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_797 (.A(n18_adj_7136), .B(n24_adj_7137), .C(n18_adj_7138), 
         .D(n4_adj_7139), .Z(n26_adj_7133)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_797.init = 16'hfffe;
    FD1P3IX reset_r_480 (.D(n29083), .SP(clk_enable_521), .CD(n29239), 
            .CK(clk), .Q(reset_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam reset_r_480.GSR = "DISABLED";
    LUT4 i8_4_lut_adj_798 (.A(\spi_data_out_r_39__N_4835[20] ), .B(n16_adj_7140), 
         .C(n17_adj_7141), .D(spi_data_out_r_39__N_4875), .Z(n22_adj_7134)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i8_4_lut_adj_798.init = 16'hfefc;
    LUT4 Select_4066_i21_2_lut (.A(\spi_data_out_r_39__N_5513[20] ), .B(spi_data_out_r_39__N_5553), 
         .Z(n21_adj_7135)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4066_i21_2_lut.init = 16'h8888;
    LUT4 Select_4066_i18_2_lut (.A(\spi_data_out_r_39__N_4496[20] ), .B(spi_data_out_r_39__N_4536), 
         .Z(n18_adj_7136)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4066_i18_2_lut.init = 16'h8888;
    LUT4 i13681_2_lut_3_lut (.A(n19439), .B(n19545), .C(n153[0]), .Z(n199[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13681_2_lut_3_lut.init = 16'h7070;
    LUT4 i10_4_lut_adj_799 (.A(\spi_data_out_r_39__N_3818[20] ), .B(n20_adj_7142), 
         .C(n5_adj_7143), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_7137)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_799.init = 16'hfefc;
    LUT4 i13898_2_lut_3_lut (.A(n19439), .B(n19545), .C(n153[1]), .Z(n199[1])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13898_2_lut_3_lut.init = 16'h7070;
    LUT4 i4_4_lut_adj_800 (.A(\spi_data_out_r_39__N_2104[20] ), .B(\spi_data_out_r_39__N_1870[20] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_7138)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_800.init = 16'heca0;
    LUT4 Select_4066_i4_2_lut (.A(\spi_data_out_r_39__N_1402[20] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_7139)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4066_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_801 (.A(\spi_data_out_r_39__N_2338[20] ), .B(\spi_data_out_r_39__N_5174[20] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_7142)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_801.init = 16'heca0;
    LUT4 Select_4066_i5_2_lut (.A(\spi_data_out_r_39__N_1636[20] ), .B(spi_data_out_r_39__N_1676), 
         .Z(n5_adj_7143)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4066_i5_2_lut.init = 16'h8888;
    LUT4 i2_4_lut_adj_802 (.A(\spi_data_out_r_39__N_934[20] ), .B(spi_data_out_r_39__N_5852[20]), 
         .C(spi_data_out_r_39__N_974), .D(spi_data_out_r_39__N_5892), .Z(n16_adj_7140)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i2_4_lut_adj_802.init = 16'heca0;
    LUT4 i13899_2_lut_3_lut (.A(n19439), .B(n19545), .C(n153[2]), .Z(n199[2])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13899_2_lut_3_lut.init = 16'h7070;
    LUT4 Select_4066_i17_2_lut (.A(\spi_data_out_r_39__N_4157[20] ), .B(spi_data_out_r_39__N_4197), 
         .Z(n17_adj_7141)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4066_i17_2_lut.init = 16'h8888;
    LUT4 i13900_2_lut_3_lut (.A(n19439), .B(n19545), .C(n153[3]), .Z(n199[3])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13900_2_lut_3_lut.init = 16'h7070;
    LUT4 i13_4_lut_adj_803 (.A(n3_adj_7144), .B(n26_adj_7145), .C(n22_adj_6773), 
         .D(n21_adj_6897), .Z(\spi_data_out_r[21] )) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i13_4_lut_adj_803.init = 16'hfffe;
    LUT4 Select_4065_i3_2_lut (.A(\spi_data_out_r_39__N_1168[21] ), .B(spi_data_out_r_39__N_1208), 
         .Z(n3_adj_7144)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4065_i3_2_lut.init = 16'h8888;
    LUT4 i12_4_lut_adj_804 (.A(n18_adj_6939), .B(n24_adj_7146), .C(n18_adj_7147), 
         .D(n4_adj_7148), .Z(n26_adj_7145)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut_adj_804.init = 16'hfffe;
    LUT4 i13901_2_lut_3_lut (.A(n19439), .B(n19545), .C(n153[4]), .Z(n199[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13901_2_lut_3_lut.init = 16'h7070;
    LUT4 i10_4_lut_adj_805 (.A(\spi_data_out_r_39__N_3818[21] ), .B(n20_adj_7149), 
         .C(n5_adj_6790), .D(spi_data_out_r_39__N_3858), .Z(n24_adj_7146)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i10_4_lut_adj_805.init = 16'hfefc;
    INV i23370 (.A(MA_Temp), .Z(MA_Temp_N_5969));
    LUT4 i13903_2_lut_3_lut (.A(n19439), .B(n19545), .C(n153[6]), .Z(n199[6])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13903_2_lut_3_lut.init = 16'h7070;
    LUT4 i13904_2_lut_3_lut (.A(n19439), .B(n19545), .C(n153[7]), .Z(n199[7])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13904_2_lut_3_lut.init = 16'h7070;
    LUT4 i4_4_lut_adj_806 (.A(\spi_data_out_r_39__N_2104[21] ), .B(\spi_data_out_r_39__N_1870[21] ), 
         .C(spi_data_out_r_39__N_2144), .D(spi_data_out_r_39__N_1910), .Z(n18_adj_7147)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i4_4_lut_adj_806.init = 16'heca0;
    LUT4 Select_4065_i4_2_lut (.A(\spi_data_out_r_39__N_1402[21] ), .B(spi_data_out_r_39__N_1442), 
         .Z(n4_adj_7148)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_4065_i4_2_lut.init = 16'h8888;
    LUT4 i6_4_lut_adj_807 (.A(\spi_data_out_r_39__N_2338[21] ), .B(\spi_data_out_r_39__N_5174[21] ), 
         .C(spi_data_out_r_39__N_2378), .D(spi_data_out_r_39__N_5214), .Z(n20_adj_7149)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i6_4_lut_adj_807.init = 16'heca0;
    
endmodule
//
// Verilog Description of module spi_slave_top
//

module spi_slave_top (spi_addr_r, clk, n29247, spi_addr, n29239, \spi_addr_r[3] , 
            \spi_addr[3] , \spi_addr_r[2] , \spi_addr[2] , \spi_addr_r[1] , 
            \spi_addr[1] , spi_cmd_r, \spi_data_r[0] , clk_enable_524, 
            n27, n29182, n13074, n29077, n29761, n27256, n29174, 
            n29211, spi_addr_valid, spi_cmd_valid, resetn_c, spi_scsn_c, 
            spi_sdo_valid_N_296, n29162, n29161, n29144, n29122, n29251, 
            n29254, n27283, n29216, n27058, n29169, n6, n13265, 
            n29214, n29127, n29118, n29130, \spi_data_r[31] , \spi_data_r[30] , 
            \spi_data_r[29] , \spi_data_r[28] , \spi_data_r[27] , \spi_data_r[26] , 
            \spi_data_r[25] , \spi_data_r[24] , \spi_data_r[23] , \spi_data_r[22] , 
            \spi_data_r[21] , \spi_data_r[20] , \spi_data_r[19] , \spi_data_r[18] , 
            \spi_data_r[17] , \spi_data_r[16] , \spi_data_r[15] , \spi_data_r[14] , 
            \spi_data_r[13] , \spi_data_r[12] , \spi_data_r[11] , \spi_data_r[10] , 
            \spi_data_r[9] , \spi_data_r[8] , \spi_data_r[7] , \spi_data_r[6] , 
            \spi_data_r[5] , \spi_data_r[4] , \spi_data_r[3] , \spi_data_r[2] , 
            \spi_data_r[1] , n27338, n29311, n27259, n29287, n29255, 
            reset_r_N_4813, clk_enable_190, n65, n29070, spi_sdo_valid_N_297, 
            \spi_data_out_r_39__N_2643[2] , n13, clear_intrpt, n4, \spi_data_out_r_39__N_934[2] , 
            n19, spi_data_out_r_39__N_974, spi_data_valid_r, spi_data_valid, 
            spi_cmd, \spi_data_out_r_39__N_4157[2] , \spi_data_out_r_39__N_1168[2] , 
            spi_data_out_r_39__N_4197, spi_data_out_r_39__N_1208, \spi_data_out_r_39__N_2927[2] , 
            \spi_data_out_r_39__N_2785[2] , clear_intrpt_adj_151, clear_intrpt_adj_152, 
            n8, n15, \spi_cmd[4] , \spi_cmd_r[6] , \spi_cmd_r[7] , 
            \spi_cmd_r[8] , \spi_cmd_r[9] , \spi_cmd_r[10] , \spi_cmd_r[11] , 
            \spi_cmd_r[12] , \spi_cmd_r[13] , \spi_cmd_r[14] , \spi_cmd_r[15] , 
            \spi_cmd[15] , \spi_data_out_r[1] , \spi_data_out_r[3] , \spi_data_out_r[4] , 
            \spi_data_out_r[5] , \spi_data_out_r[6] , \spi_data_out_r[7] , 
            \spi_data_out_r[8] , \spi_data_out_r[9] , \spi_data_out_r[10] , 
            \spi_data_out_r[11] , \spi_data_out_r[12] , \spi_data_out_r[13] , 
            \spi_data_out_r[14] , \spi_data_out_r[15] , \spi_data_out_r[16] , 
            \spi_data_out_r[17] , \spi_data_out_r[18] , \spi_data_out_r[19] , 
            \spi_data_out_r[20] , \spi_data_out_r[21] , \spi_data_out_r[22] , 
            \spi_data_out_r[23] , \spi_data_out_r[24] , \spi_data_out_r[25] , 
            \spi_data_out_r[26] , \spi_data_out_r[27] , \spi_data_out_r[28] , 
            \spi_data_out_r[29] , \spi_data_out_r[30] , \spi_data_out_r[31] , 
            \spi_data_out_r[32] , \spi_data_out_r[33] , \spi_data_out_r[34] , 
            \spi_data_out_r[35] , \spi_data_out_r[36] , \spi_data_out_r[37] , 
            \spi_data_out_r[38] , \spi_data_out_r[39] , \spi_data_out_r_39__N_5174[2] , 
            \spi_data_out_r_39__N_3818[2] , spi_data_out_r_39__N_5214, spi_data_out_r_39__N_3858, 
            \spi_data_out_r_39__N_5852[2] , n11, spi_data_out_r_39__N_5892, 
            \spi_data_out_r_39__N_4496[2] , \spi_data_out_r_39__N_1870[2] , 
            spi_data_out_r_39__N_4536, spi_data_out_r_39__N_1910, \spi_data_out_r_39__N_5513[2] , 
            \spi_data_out_r_39__N_1636[2] , spi_data_out_r_39__N_5553, spi_data_out_r_39__N_1676, 
            \spi_data_out_r_39__N_2104[2] , \spi_data_out_r_39__N_2572[2] , 
            spi_data_out_r_39__N_2144, clear_intrpt_adj_153, n29075, n29078, 
            n29079, n29080, n27286, n65_adj_154, n29092, \spi_data_out_r_39__N_2927[0] , 
            n17, n3, n20, \spi_data_out_r_39__N_3818[0] , n4_adj_155, 
            \spi_data_out_r_39__N_1870[0] , \spi_data_out_r_39__N_2785[0] , 
            n15_adj_156, n2, \spi_data_out_r_39__N_4496[0] , n11_adj_157, 
            \spi_data_out_r_39__N_4835[0] , n21, spi_data_out_r_39__N_4875, 
            \spi_data_out_r_39__N_770[0] , \spi_data_out_r_39__N_5852[0] , 
            spi_data_out_r_39__N_810, \spi_data_out_r_39__N_2338[0] , \spi_data_out_r_39__N_2572[0] , 
            spi_data_out_r_39__N_2378, \spi_data_out_r_39__N_2104[0] , \spi_data_out_r_39__N_2856[0] , 
            clear_intrpt_adj_158, \spi_data_out_r_39__N_1636[0] , \spi_data_out_r_39__N_2643[0] , 
            n29089, clk_enable_206, n29096, n29213, n29097, n29106, 
            n29123, n29762, n29757, GND_net, spi_mosi_oe, spi_mosi_o, 
            spi_miso_oe, spi_miso_o, spi_clk_oe, spi_clk_o, spi_mosi_i, 
            spi_miso_i, spi_clk_i, VCC_net, mem_rdata_update_N_729, 
            quad_set_complete, clk_enable_518, n27225, clk_enable_398, 
            n29102, clk_enable_188, clk_enable_303, n32, \quad_homing[1] , 
            n27657, n24, clk_enable_179, clk_enable_182, intrpt_out_N_2848, 
            n29100, clk_enable_185, n29134, clk_enable_509, EM_STOP, 
            clk_enable_306, n29101, clk_enable_186, quad_set_complete_adj_159, 
            n29120, clk_enable_505, clk_enable_76, n29104, clk_enable_436, 
            n19233, clk_enable_184, clk_enable_204, intrpt_out_N_2635, 
            n29288, clk_enable_183, clk_enable_271, n29083, clk_enable_521, 
            quad_set_valid, n66, n21446, clk_1MHz_enable_171, n29124, 
            clk_enable_197, n26948, n13_adj_160, n12714, n27301, clk_enable_193, 
            clk_enable_200, n29307, clk_enable_499, n27240, clk_enable_32, 
            quad_set_complete_adj_161, clk_enable_520, n29286, clk_enable_77, 
            intrpt_out_N_2706, quad_set_valid_adj_162, n79, n20819, 
            clk_1MHz_enable_340, n27285, n29110, clk_enable_340, n31, 
            \quad_homing[1]_adj_163 , n5, n26, n27234, clk_enable_174, 
            clk_enable_171, clk_enable_172, clk_enable_435, n29082, 
            clk_enable_506, clk_enable_269, clk_enable_167, clk_enable_28, 
            clk_enable_131, intrpt_out_N_2919, clk_enable_194, clk_enable_177, 
            clk_enable_189, clk_enable_180, clk_enable_162, clk_enable_166, 
            n29256, clk_enable_175, clk_enable_176, quad_set_complete_adj_164, 
            n29105, clk_enable_502, clk_enable_526, clk_enable_342, 
            clk_enable_202, intrpt_out_N_2990, clk_enable_201, clk_enable_467, 
            clk_enable_191, clk_enable_187, clk_enable_192, quad_set_complete_adj_165, 
            clk_enable_519, clk_enable_170, clk_enable_286, clk_enable_359, 
            reset_r_N_4474, clk_enable_307, clear_intrpt_adj_166, intrpt_out_N_3061, 
            clk_enable_86, clk_enable_181, clk_enable_288, clk_enable_433, 
            clk_enable_434, quad_set_complete_adj_167, clk_enable_501, 
            n29205, clk_enable_169, clear_intrpt_adj_168, intrpt_out_N_2777, 
            clk_enable_400, clk_enable_402, quad_set_complete_adj_169, 
            clk_enable_503, clk_enable_30, n9633, n27465, n26928, 
            n29141, n29126, n27618, n29114, clk_enable_20, \spi_cmd[0] , 
            n31_adj_170) /* synthesis syn_module_defined=1 */ ;
    output [7:0]spi_addr_r;
    input clk;
    output n29247;
    output [7:0]spi_addr;
    output n29239;
    output \spi_addr_r[3] ;
    output \spi_addr[3] ;
    output \spi_addr_r[2] ;
    output \spi_addr[2] ;
    output \spi_addr_r[1] ;
    output \spi_addr[1] ;
    output [15:0]spi_cmd_r;
    output \spi_data_r[0] ;
    input clk_enable_524;
    output n27;
    output n29182;
    input n13074;
    output n29077;
    output n29761;
    output n27256;
    output n29174;
    output n29211;
    output spi_addr_valid;
    output spi_cmd_valid;
    input resetn_c;
    input spi_scsn_c;
    output spi_sdo_valid_N_296;
    output n29162;
    input n29161;
    output n29144;
    output n29122;
    output n29251;
    output n29254;
    output n27283;
    output n29216;
    input n27058;
    input n29169;
    output n6;
    input n13265;
    input n29214;
    output n29127;
    output n29118;
    output n29130;
    output \spi_data_r[31] ;
    output \spi_data_r[30] ;
    output \spi_data_r[29] ;
    output \spi_data_r[28] ;
    output \spi_data_r[27] ;
    output \spi_data_r[26] ;
    output \spi_data_r[25] ;
    output \spi_data_r[24] ;
    output \spi_data_r[23] ;
    output \spi_data_r[22] ;
    output \spi_data_r[21] ;
    output \spi_data_r[20] ;
    output \spi_data_r[19] ;
    output \spi_data_r[18] ;
    output \spi_data_r[17] ;
    output \spi_data_r[16] ;
    output \spi_data_r[15] ;
    output \spi_data_r[14] ;
    output \spi_data_r[13] ;
    output \spi_data_r[12] ;
    output \spi_data_r[11] ;
    output \spi_data_r[10] ;
    output \spi_data_r[9] ;
    output \spi_data_r[8] ;
    output \spi_data_r[7] ;
    output \spi_data_r[6] ;
    output \spi_data_r[5] ;
    output \spi_data_r[4] ;
    output \spi_data_r[3] ;
    output \spi_data_r[2] ;
    output \spi_data_r[1] ;
    output n27338;
    output n29311;
    output n27259;
    input n29287;
    input n29255;
    input reset_r_N_4813;
    output clk_enable_190;
    input n65;
    output n29070;
    input spi_sdo_valid_N_297;
    input \spi_data_out_r_39__N_2643[2] ;
    input n13;
    input clear_intrpt;
    input n4;
    input \spi_data_out_r_39__N_934[2] ;
    input n19;
    input spi_data_out_r_39__N_974;
    output spi_data_valid_r;
    output spi_data_valid;
    output [15:0]spi_cmd;
    input \spi_data_out_r_39__N_4157[2] ;
    input \spi_data_out_r_39__N_1168[2] ;
    input spi_data_out_r_39__N_4197;
    input spi_data_out_r_39__N_1208;
    input \spi_data_out_r_39__N_2927[2] ;
    input \spi_data_out_r_39__N_2785[2] ;
    input clear_intrpt_adj_151;
    input clear_intrpt_adj_152;
    input n8;
    input n15;
    output \spi_cmd[4] ;
    output \spi_cmd_r[6] ;
    output \spi_cmd_r[7] ;
    output \spi_cmd_r[8] ;
    output \spi_cmd_r[9] ;
    output \spi_cmd_r[10] ;
    output \spi_cmd_r[11] ;
    output \spi_cmd_r[12] ;
    output \spi_cmd_r[13] ;
    output \spi_cmd_r[14] ;
    output \spi_cmd_r[15] ;
    output \spi_cmd[15] ;
    input \spi_data_out_r[1] ;
    input \spi_data_out_r[3] ;
    input \spi_data_out_r[4] ;
    input \spi_data_out_r[5] ;
    input \spi_data_out_r[6] ;
    input \spi_data_out_r[7] ;
    input \spi_data_out_r[8] ;
    input \spi_data_out_r[9] ;
    input \spi_data_out_r[10] ;
    input \spi_data_out_r[11] ;
    input \spi_data_out_r[12] ;
    input \spi_data_out_r[13] ;
    input \spi_data_out_r[14] ;
    input \spi_data_out_r[15] ;
    input \spi_data_out_r[16] ;
    input \spi_data_out_r[17] ;
    input \spi_data_out_r[18] ;
    input \spi_data_out_r[19] ;
    input \spi_data_out_r[20] ;
    input \spi_data_out_r[21] ;
    input \spi_data_out_r[22] ;
    input \spi_data_out_r[23] ;
    input \spi_data_out_r[24] ;
    input \spi_data_out_r[25] ;
    input \spi_data_out_r[26] ;
    input \spi_data_out_r[27] ;
    input \spi_data_out_r[28] ;
    input \spi_data_out_r[29] ;
    input \spi_data_out_r[30] ;
    input \spi_data_out_r[31] ;
    input \spi_data_out_r[32] ;
    input \spi_data_out_r[33] ;
    input \spi_data_out_r[34] ;
    input \spi_data_out_r[35] ;
    input \spi_data_out_r[36] ;
    input \spi_data_out_r[37] ;
    input \spi_data_out_r[38] ;
    input \spi_data_out_r[39] ;
    input \spi_data_out_r_39__N_5174[2] ;
    input \spi_data_out_r_39__N_3818[2] ;
    input spi_data_out_r_39__N_5214;
    input spi_data_out_r_39__N_3858;
    input \spi_data_out_r_39__N_5852[2] ;
    input n11;
    input spi_data_out_r_39__N_5892;
    input \spi_data_out_r_39__N_4496[2] ;
    input \spi_data_out_r_39__N_1870[2] ;
    input spi_data_out_r_39__N_4536;
    input spi_data_out_r_39__N_1910;
    input \spi_data_out_r_39__N_5513[2] ;
    input \spi_data_out_r_39__N_1636[2] ;
    input spi_data_out_r_39__N_5553;
    input spi_data_out_r_39__N_1676;
    input \spi_data_out_r_39__N_2104[2] ;
    input \spi_data_out_r_39__N_2572[2] ;
    input spi_data_out_r_39__N_2144;
    input clear_intrpt_adj_153;
    output n29075;
    output n29078;
    output n29079;
    output n29080;
    input n27286;
    input n65_adj_154;
    output n29092;
    input \spi_data_out_r_39__N_2927[0] ;
    input n17;
    input n3;
    input n20;
    input \spi_data_out_r_39__N_3818[0] ;
    input n4_adj_155;
    input \spi_data_out_r_39__N_1870[0] ;
    input \spi_data_out_r_39__N_2785[0] ;
    input n15_adj_156;
    input n2;
    input \spi_data_out_r_39__N_4496[0] ;
    input n11_adj_157;
    input \spi_data_out_r_39__N_4835[0] ;
    input n21;
    input spi_data_out_r_39__N_4875;
    input \spi_data_out_r_39__N_770[0] ;
    input \spi_data_out_r_39__N_5852[0] ;
    input spi_data_out_r_39__N_810;
    input \spi_data_out_r_39__N_2338[0] ;
    input \spi_data_out_r_39__N_2572[0] ;
    input spi_data_out_r_39__N_2378;
    input \spi_data_out_r_39__N_2104[0] ;
    input \spi_data_out_r_39__N_2856[0] ;
    input clear_intrpt_adj_158;
    input \spi_data_out_r_39__N_1636[0] ;
    input \spi_data_out_r_39__N_2643[0] ;
    output n29089;
    output clk_enable_206;
    output n29096;
    input n29213;
    output n29097;
    output n29106;
    output n29123;
    output n29762;
    input n29757;
    input GND_net;
    output spi_mosi_oe;
    output spi_mosi_o;
    output spi_miso_oe;
    output spi_miso_o;
    output spi_clk_oe;
    output spi_clk_o;
    input spi_mosi_i;
    input spi_miso_i;
    input spi_clk_i;
    input VCC_net;
    output mem_rdata_update_N_729;
    input quad_set_complete;
    output clk_enable_518;
    input n27225;
    output clk_enable_398;
    input n29102;
    output clk_enable_188;
    output clk_enable_303;
    input n32;
    input \quad_homing[1] ;
    input n27657;
    output n24;
    output clk_enable_179;
    output clk_enable_182;
    output intrpt_out_N_2848;
    input n29100;
    output clk_enable_185;
    input n29134;
    output clk_enable_509;
    input EM_STOP;
    output clk_enable_306;
    input n29101;
    output clk_enable_186;
    input quad_set_complete_adj_159;
    input n29120;
    output clk_enable_505;
    output clk_enable_76;
    input n29104;
    output clk_enable_436;
    input n19233;
    output clk_enable_184;
    output clk_enable_204;
    output intrpt_out_N_2635;
    input n29288;
    output clk_enable_183;
    output clk_enable_271;
    input n29083;
    output clk_enable_521;
    input quad_set_valid;
    input n66;
    input n21446;
    output clk_1MHz_enable_171;
    input n29124;
    output clk_enable_197;
    input n26948;
    input n13_adj_160;
    input n12714;
    output n27301;
    output clk_enable_193;
    output clk_enable_200;
    input n29307;
    output clk_enable_499;
    input n27240;
    output clk_enable_32;
    input quad_set_complete_adj_161;
    output clk_enable_520;
    input n29286;
    output clk_enable_77;
    output intrpt_out_N_2706;
    input quad_set_valid_adj_162;
    input n79;
    input n20819;
    output clk_1MHz_enable_340;
    input n27285;
    input n29110;
    output clk_enable_340;
    input n31;
    input \quad_homing[1]_adj_163 ;
    input n5;
    output n26;
    input n27234;
    output clk_enable_174;
    output clk_enable_171;
    output clk_enable_172;
    output clk_enable_435;
    input n29082;
    output clk_enable_506;
    output clk_enable_269;
    output clk_enable_167;
    output clk_enable_28;
    output clk_enable_131;
    output intrpt_out_N_2919;
    output clk_enable_194;
    output clk_enable_177;
    output clk_enable_189;
    output clk_enable_180;
    output clk_enable_162;
    output clk_enable_166;
    input n29256;
    output clk_enable_175;
    output clk_enable_176;
    input quad_set_complete_adj_164;
    input n29105;
    output clk_enable_502;
    output clk_enable_526;
    output clk_enable_342;
    output clk_enable_202;
    output intrpt_out_N_2990;
    output clk_enable_201;
    output clk_enable_467;
    output clk_enable_191;
    output clk_enable_187;
    output clk_enable_192;
    input quad_set_complete_adj_165;
    output clk_enable_519;
    output clk_enable_170;
    output clk_enable_286;
    output clk_enable_359;
    input reset_r_N_4474;
    output clk_enable_307;
    input clear_intrpt_adj_166;
    output intrpt_out_N_3061;
    output clk_enable_86;
    output clk_enable_181;
    output clk_enable_288;
    output clk_enable_433;
    output clk_enable_434;
    input quad_set_complete_adj_167;
    output clk_enable_501;
    input n29205;
    output clk_enable_169;
    input clear_intrpt_adj_168;
    output intrpt_out_N_2777;
    output clk_enable_400;
    output clk_enable_402;
    input quad_set_complete_adj_169;
    output clk_enable_503;
    output clk_enable_30;
    input n9633;
    output n27465;
    output n26928;
    output n29141;
    output n29126;
    output n27618;
    input n29114;
    output clk_enable_20;
    output \spi_cmd[0] ;
    output n31_adj_170;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire spi_clk_i /* synthesis is_clock=1 */ ;   // c:/s_links/sources/config_mcm/ip/spi_slave_efb.v(34[10:19])
    
    wire clk_enable_14;
    wire [39:0]spi_sdo_r;   // c:/s_links/sources/spi_slave_top.v(66[23:32])
    
    wire clk_enable_523, n27177;
    wire [7:0]spi_addr_r_c;   // c:/s_links/sources/mcm_top.v(84[28:38])
    wire [7:0]spi_addr_c;   // c:/s_links/sources/mcm_top.v(89[28:36])
    wire [39:0]spi_sdo;   // c:/s_links/sources/spi_slave_top.v(74[23:30])
    
    wire clk_enable_305;
    wire [39:0]spi_sdo_39__N_145;
    
    wire spi_sdo_valid;
    wire [39:0]mem_rdata_7__N_185;
    
    wire n4_c;
    wire [39:0]spi_data;   // c:/s_links/sources/spi_slave_top.v(70[23:31])
    
    wire n27176, n29107, clk_enable_357, n29069, n29242, n27201, 
        n29175, n27243, clk_enable_341, spi_scsn_dly, clk_enable_196;
    wire [15:0]spi_cmd_r_c;   // c:/s_links/sources/mcm_top.v(83[27:36])
    
    wire spi_addr_valid_r_N_303, n27280, n29119, n29129, n29121, n29081, 
        n29095, n27178, n27172, n27179, n27173, n27174, n27175;
    wire [7:0]mem_rdata;   // c:/s_links/sources/spi_slave_top.v(64[32:41])
    
    wire n35, n40, n36, n28, n31_c, n38, n22, n30, n34, n24_c;
    wire [15:0]spi_cmd_c;   // c:/s_links/sources/mcm_top.v(88[27:34])
    
    wire n10988, n26_c, n29074, n29072, n29071, n37, n42, n38_adj_6731, 
        n30_adj_6732, n40_adj_6733, n34_adj_6734, n32_c, n36_adj_6737, 
        n26_adj_6738, n24_adj_6739, n28_adj_6741, n60, n29086, n29090, 
        n29111, wb_cyc_i, clk_enable_95, wb_cyc_i_N_339;
    wire [7:0]wb_adr_i;   // c:/s_links/sources/spi_slave_top.v(47[44:52])
    wire [7:0]address;   // c:/s_links/sources/spi_slave_top.v(52[44:51])
    
    wire wb_we_i, wb_we_i_N_344;
    wire [7:0]wb_dat_i;   // c:/s_links/sources/spi_slave_top.v(48[44:52])
    wire [7:0]wr_data;   // c:/s_links/sources/spi_slave_top.v(54[44:51])
    
    wire wb_sm, n28767, n29268;
    wire [7:0]address_7__N_549;
    
    wire spi_cmd_start;
    wire [7:0]address_7__N_565;
    
    wire wr_en, wr_en_N_355;
    wire [7:0]wb_dat_o;   // c:/s_links/sources/spi_slave_top.v(49[44:52])
    wire [15:0]n2713;
    
    wire spi_addr_valid_N_732, n29176, n29179, n7083, clk_enable_309, 
        clk_enable_516;
    
    FD1P3IX spi_addr_r__i0 (.D(spi_addr[0]), .SP(clk_enable_14), .CD(n29247), 
            .CK(clk), .Q(spi_addr_r[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i0.GSR = "DISABLED";
    FD1P3AX spi_sdo_r__i1 (.D(n27177), .SP(clk_enable_523), .CK(clk), 
            .Q(spi_sdo_r[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i1.GSR = "DISABLED";
    FD1P3IX spi_addr_r__i7 (.D(spi_addr_c[7]), .SP(clk_enable_14), .CD(n29247), 
            .CK(clk), .Q(spi_addr_r_c[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i7.GSR = "DISABLED";
    FD1P3IX spi_addr_r__i6 (.D(spi_addr_c[6]), .SP(clk_enable_14), .CD(n29247), 
            .CK(clk), .Q(spi_addr_r_c[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i6.GSR = "DISABLED";
    FD1P3IX spi_sdo__i2 (.D(spi_sdo_39__N_145[2]), .SP(clk_enable_305), 
            .CD(n29239), .CK(clk), .Q(spi_sdo[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i2.GSR = "DISABLED";
    FD1P3IX spi_addr_r__i5 (.D(spi_addr_c[5]), .SP(clk_enable_14), .CD(n29247), 
            .CK(clk), .Q(spi_addr_r_c[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i5.GSR = "DISABLED";
    FD1P3IX spi_addr_r__i4 (.D(spi_addr_c[4]), .SP(clk_enable_14), .CD(n29247), 
            .CK(clk), .Q(spi_addr_r_c[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i4.GSR = "DISABLED";
    FD1P3IX spi_addr_r__i3 (.D(\spi_addr[3] ), .SP(clk_enable_14), .CD(n29247), 
            .CK(clk), .Q(\spi_addr_r[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i3.GSR = "DISABLED";
    FD1P3IX spi_addr_r__i2 (.D(\spi_addr[2] ), .SP(clk_enable_14), .CD(n29247), 
            .CK(clk), .Q(\spi_addr_r[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i2.GSR = "DISABLED";
    FD1P3IX spi_addr_r__i1 (.D(\spi_addr[1] ), .SP(clk_enable_14), .CD(n29247), 
            .CK(clk), .Q(\spi_addr_r[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_r__i1.GSR = "DISABLED";
    LUT4 mux_18_i17_3_lut (.A(spi_sdo_r[8]), .B(spi_sdo[16]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i17_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(spi_cmd_r[2]), .B(\spi_addr_r[2] ), .Z(n4_c)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut.init = 16'h8888;
    FD1P3IX spi_data_r__i0 (.D(spi_data[0]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i0.GSR = "DISABLED";
    LUT4 i3_4_lut (.A(spi_addr_r_c[7]), .B(spi_addr_r_c[5]), .C(spi_addr_r_c[6]), 
         .D(spi_addr_r_c[4]), .Z(n27)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    FD1P3IX spi_sdo_r__i17 (.D(mem_rdata_7__N_185[17]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i17.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i16 (.D(mem_rdata_7__N_185[16]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i16.GSR = "DISABLED";
    FD1P3AX spi_sdo_r__i2 (.D(n27176), .SP(clk_enable_523), .CK(clk), 
            .Q(spi_sdo_r[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i2.GSR = "DISABLED";
    LUT4 i2_3_lut_rep_349_4_lut (.A(spi_cmd_r[2]), .B(n29107), .C(n29182), 
         .D(n13074), .Z(n29077)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i2_3_lut_rep_349_4_lut.init = 16'h0400;
    FD1P3IX spi_cmd_r__i0 (.D(n29761), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(spi_cmd_r[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i0.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i15 (.D(mem_rdata_7__N_185[15]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i15.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_341_3_lut_4_lut (.A(spi_cmd_r[2]), .B(n29107), .C(n27256), 
         .D(n29174), .Z(n29069)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_341_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_rep_514 (.A(spi_cmd_r[1]), .B(spi_addr_r[0]), .Z(n29242)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_514.init = 16'h8888;
    LUT4 i1_2_lut_rep_483_3_lut (.A(spi_cmd_r[1]), .B(spi_addr_r[0]), .C(spi_cmd_r[0]), 
         .Z(n29211)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_483_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_3_lut (.A(spi_cmd_r[1]), .B(spi_addr_r[0]), .C(spi_cmd_r[3]), 
         .Z(n27256)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut (.A(spi_cmd_r[1]), .B(spi_addr_r[0]), .C(\spi_addr_r[1] ), 
         .D(spi_cmd_r[3]), .Z(n27201)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_rep_447_3_lut (.A(spi_cmd_r[1]), .B(spi_addr_r[0]), .C(spi_cmd_r[3]), 
         .Z(n29175)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_447_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_3_lut_4_lut_adj_553 (.A(spi_cmd_r[1]), .B(spi_addr_r[0]), 
         .C(\spi_addr_r[1] ), .D(spi_cmd_r[3]), .Z(n27243)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_3_lut_4_lut_adj_553.init = 16'h0080;
    LUT4 i22876_2_lut_rep_518 (.A(spi_addr_valid), .B(spi_cmd_valid), .Z(clk_enable_341)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/spi_slave_top.v(137[8] 149[6])
    defparam i22876_2_lut_rep_518.init = 16'hdddd;
    LUT4 i2728_2_lut_2_lut_3_lut (.A(spi_addr_valid), .B(spi_cmd_valid), 
         .C(n29247), .Z(clk_enable_14)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // c:/s_links/sources/spi_slave_top.v(137[8] 149[6])
    defparam i2728_2_lut_2_lut_3_lut.init = 16'hf2f2;
    LUT4 wb_rst_i_I_0_3_lut_rep_519 (.A(resetn_c), .B(spi_scsn_c), .C(spi_scsn_dly), 
         .Z(n29247)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(124[7:26])
    defparam wb_rst_i_I_0_3_lut_rep_519.init = 16'h5d5d;
    LUT4 i2730_2_lut_4_lut (.A(resetn_c), .B(spi_scsn_c), .C(spi_scsn_dly), 
         .D(spi_cmd_valid), .Z(clk_enable_196)) /* synthesis lut_function=(!(A (B (C (D))+!B (D)))) */ ;   // c:/s_links/sources/spi_slave_top.v(124[7:26])
    defparam i2730_2_lut_4_lut.init = 16'h5dff;
    LUT4 i2727_2_lut_4_lut (.A(resetn_c), .B(spi_scsn_c), .C(spi_scsn_dly), 
         .D(spi_cmd_valid), .Z(clk_enable_357)) /* synthesis lut_function=((B ((D)+!C)+!B (D))+!A) */ ;   // c:/s_links/sources/spi_slave_top.v(124[7:26])
    defparam i2727_2_lut_4_lut.init = 16'hff5d;
    FD1S3IX spi_sdo_valid_52 (.D(spi_sdo_valid_N_296), .CK(clk), .CD(n29239), 
            .Q(spi_sdo_valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo_valid_52.GSR = "DISABLED";
    FD1S3IX spi_scsn_dly_59 (.D(spi_scsn_c), .CK(clk), .CD(n29239), .Q(spi_scsn_dly)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(153[9] 158[5])
    defparam spi_scsn_dly_59.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_394_3_lut_4_lut (.A(n29162), .B(n29161), .C(n29144), 
         .D(spi_cmd_r[2]), .Z(n29122)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_394_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_523 (.A(spi_cmd_r_c[5]), .B(spi_cmd_r_c[4]), .Z(n29251)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_523.init = 16'heeee;
    LUT4 i13636_2_lut_rep_454_3_lut (.A(spi_cmd_r_c[5]), .B(spi_cmd_r_c[4]), 
         .C(spi_cmd_r[3]), .Z(n29182)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i13636_2_lut_rep_454_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_526 (.A(spi_cmd_r[3]), .B(\spi_addr_r[1] ), .Z(n29254)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_526.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_554 (.A(spi_cmd_r[3]), .B(\spi_addr_r[1] ), 
         .C(spi_addr_r[0]), .D(spi_cmd_r[1]), .Z(n27283)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_3_lut_4_lut_adj_554.init = 16'h8000;
    FD1P3IX spi_addr_valid_r_56 (.D(spi_addr_valid_r_N_303), .SP(clk_enable_196), 
            .CD(n29247), .CK(clk), .Q(spi_sdo_valid_N_296)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_addr_valid_r_56.GSR = "DISABLED";
    LUT4 i3_4_lut_adj_555 (.A(n29216), .B(n27058), .C(n29169), .D(n27280), 
         .Z(n6)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i3_4_lut_adj_555.init = 16'h0800;
    LUT4 i1_2_lut_rep_416 (.A(\spi_addr_r[3] ), .B(n13265), .Z(n29144)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_416.init = 16'h4444;
    LUT4 i1_2_lut_rep_391_3_lut_4_lut (.A(\spi_addr_r[3] ), .B(n13265), 
         .C(n29214), .D(spi_cmd_r[2]), .Z(n29119)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_391_3_lut_4_lut.init = 16'h0004;
    LUT4 i1_2_lut_rep_399_3_lut (.A(\spi_addr_r[3] ), .B(n13265), .C(spi_cmd_r[2]), 
         .Z(n29127)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_399_3_lut.init = 16'h0404;
    LUT4 i1_2_lut_rep_390_3_lut_4_lut (.A(\spi_addr_r[3] ), .B(n13265), 
         .C(n29174), .D(spi_cmd_r[2]), .Z(n29118)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_390_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_401_3_lut (.A(\spi_addr_r[3] ), .B(n13265), .C(spi_cmd_r[2]), 
         .Z(n29129)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_401_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_402_3_lut (.A(\spi_addr_r[3] ), .B(n13265), .C(n27), 
         .Z(n29130)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_402_3_lut.init = 16'h0404;
    LUT4 i1_2_lut_rep_393_3_lut_4_lut (.A(\spi_addr_r[3] ), .B(n13265), 
         .C(\spi_addr_r[2] ), .D(n27), .Z(n29121)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_393_3_lut_4_lut.init = 16'h0040;
    FD1P3IX spi_data_r__i31 (.D(spi_data[31]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i31.GSR = "DISABLED";
    FD1P3IX spi_data_r__i30 (.D(spi_data[30]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i30.GSR = "DISABLED";
    FD1P3IX spi_data_r__i29 (.D(spi_data[29]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i29.GSR = "DISABLED";
    FD1P3IX spi_data_r__i28 (.D(spi_data[28]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i28.GSR = "DISABLED";
    FD1P3IX spi_data_r__i27 (.D(spi_data[27]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i27.GSR = "DISABLED";
    FD1P3IX spi_data_r__i26 (.D(spi_data[26]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i26.GSR = "DISABLED";
    FD1P3IX spi_data_r__i25 (.D(spi_data[25]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i25.GSR = "DISABLED";
    FD1P3IX spi_data_r__i24 (.D(spi_data[24]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i24.GSR = "DISABLED";
    FD1P3IX spi_data_r__i23 (.D(spi_data[23]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i23.GSR = "DISABLED";
    FD1P3IX spi_data_r__i22 (.D(spi_data[22]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i22.GSR = "DISABLED";
    FD1P3IX spi_data_r__i21 (.D(spi_data[21]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i21.GSR = "DISABLED";
    FD1P3IX spi_data_r__i20 (.D(spi_data[20]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i20.GSR = "DISABLED";
    FD1P3IX spi_data_r__i19 (.D(spi_data[19]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i19.GSR = "DISABLED";
    FD1P3IX spi_data_r__i18 (.D(spi_data[18]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i18.GSR = "DISABLED";
    FD1P3IX spi_data_r__i17 (.D(spi_data[17]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i17.GSR = "DISABLED";
    FD1P3IX spi_data_r__i16 (.D(spi_data[16]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i16.GSR = "DISABLED";
    FD1P3IX spi_data_r__i15 (.D(spi_data[15]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i15.GSR = "DISABLED";
    FD1P3IX spi_data_r__i14 (.D(spi_data[14]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i14.GSR = "DISABLED";
    FD1P3IX spi_data_r__i13 (.D(spi_data[13]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i13.GSR = "DISABLED";
    FD1P3IX spi_data_r__i12 (.D(spi_data[12]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i12.GSR = "DISABLED";
    FD1P3IX spi_data_r__i11 (.D(spi_data[11]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i11.GSR = "DISABLED";
    FD1P3IX spi_data_r__i10 (.D(spi_data[10]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i10.GSR = "DISABLED";
    FD1P3IX spi_data_r__i9 (.D(spi_data[9]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i9.GSR = "DISABLED";
    FD1P3IX spi_data_r__i8 (.D(spi_data[8]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i8.GSR = "DISABLED";
    FD1P3IX spi_data_r__i7 (.D(spi_data[7]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i7.GSR = "DISABLED";
    FD1P3IX spi_data_r__i6 (.D(spi_data[6]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i6.GSR = "DISABLED";
    FD1P3IX spi_data_r__i5 (.D(spi_data[5]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i5.GSR = "DISABLED";
    FD1P3IX spi_data_r__i4 (.D(spi_data[4]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i4.GSR = "DISABLED";
    FD1P3IX spi_data_r__i3 (.D(spi_data[3]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i3.GSR = "DISABLED";
    FD1P3IX spi_data_r__i2 (.D(spi_data[2]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i2.GSR = "DISABLED";
    FD1P3IX spi_data_r__i1 (.D(spi_data[1]), .SP(clk_enable_524), .CD(n29247), 
            .CK(clk), .Q(\spi_data_r[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i1.GSR = "DISABLED";
    LUT4 i1_2_lut_adj_556 (.A(\spi_addr_r[3] ), .B(n13265), .Z(n27280)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_adj_556.init = 16'h8888;
    LUT4 i2_3_lut_4_lut (.A(n29182), .B(n29107), .C(resetn_c), .D(spi_cmd_r[2]), 
         .Z(n27338)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i2_3_lut_4_lut.init = 16'hffbf;
    LUT4 mux_18_i18_3_lut (.A(spi_sdo_r[9]), .B(spi_sdo[17]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i18_3_lut.init = 16'hcaca;
    LUT4 mux_18_i16_3_lut (.A(spi_sdo_r[7]), .B(spi_sdo[15]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i16_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut_adj_557 (.A(spi_cmd_r[3]), .B(n29311), .C(n29242), 
         .D(spi_cmd_r[0]), .Z(n27259)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_3_lut_4_lut_adj_557.init = 16'h0040;
    LUT4 i1_2_lut_rep_434_3_lut_4_lut (.A(spi_cmd_r[3]), .B(n29311), .C(spi_cmd_r[0]), 
         .D(n29287), .Z(n29162)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_434_3_lut_4_lut.init = 16'h0400;
    LUT4 i4786_3_lut_4_lut (.A(n29255), .B(n29081), .C(resetn_c), .D(reset_r_N_4813), 
         .Z(clk_enable_190)) /* synthesis lut_function=(A (D)+!A !(B (C+!(D))+!B !(D))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i4786_3_lut_4_lut.init = 16'hbf00;
    LUT4 i1_2_lut_rep_367 (.A(n65), .B(\spi_addr_r[2] ), .Z(n29095)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_367.init = 16'h2222;
    LUT4 i1_2_lut_rep_353_3_lut (.A(n65), .B(\spi_addr_r[2] ), .C(spi_cmd_r[2]), 
         .Z(n29081)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_353_3_lut.init = 16'h0202;
    LUT4 i1_2_lut_rep_342_3_lut_4_lut (.A(n65), .B(\spi_addr_r[2] ), .C(n29255), 
         .D(spi_cmd_r[2]), .Z(n29070)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_342_3_lut_4_lut.init = 16'h0002;
    FD1P3IX spi_sdo_r__i14 (.D(mem_rdata_7__N_185[14]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i14.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_558 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[1]), 
         .Z(n27177)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_558.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_559 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[2]), 
         .Z(n27176)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_559.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_560 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[0]), 
         .Z(n27178)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_560.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_561 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[7]), 
         .Z(n27172)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_561.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_562 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[6]), 
         .Z(n27179)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_562.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_563 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[5]), 
         .Z(n27173)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_563.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_564 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[4]), 
         .Z(n27174)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_564.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_565 (.A(resetn_c), .B(spi_sdo_valid), .C(spi_sdo[3]), 
         .Z(n27175)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_565.init = 16'h8080;
    FD1P3AX spi_sdo_r__i0 (.D(n27178), .SP(clk_enable_523), .CK(clk), 
            .Q(spi_sdo_r[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i0.GSR = "DISABLED";
    FD1P3IX spi_sdo__i0 (.D(spi_sdo_39__N_145[0]), .SP(clk_enable_305), 
            .CD(n29239), .CK(clk), .Q(spi_sdo[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i0.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i39 (.D(mem_rdata_7__N_185[39]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(mem_rdata[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i39.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i38 (.D(mem_rdata_7__N_185[38]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(mem_rdata[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i38.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i37 (.D(mem_rdata_7__N_185[37]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(mem_rdata[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i37.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i36 (.D(mem_rdata_7__N_185[36]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(mem_rdata[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i36.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i35 (.D(mem_rdata_7__N_185[35]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(mem_rdata[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i35.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i34 (.D(mem_rdata_7__N_185[34]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(mem_rdata[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i34.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i33 (.D(mem_rdata_7__N_185[33]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(mem_rdata[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i33.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i32 (.D(mem_rdata_7__N_185[32]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(mem_rdata[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i32.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i31 (.D(mem_rdata_7__N_185[31]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i31.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i30 (.D(mem_rdata_7__N_185[30]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i30.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i29 (.D(mem_rdata_7__N_185[29]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i29.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i28 (.D(mem_rdata_7__N_185[28]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i28.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i27 (.D(mem_rdata_7__N_185[27]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i27.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i26 (.D(mem_rdata_7__N_185[26]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i26.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i25 (.D(mem_rdata_7__N_185[25]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i25.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i24 (.D(mem_rdata_7__N_185[24]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i24.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i23 (.D(mem_rdata_7__N_185[23]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i23.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i22 (.D(mem_rdata_7__N_185[22]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i22.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i21 (.D(mem_rdata_7__N_185[21]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i21.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i20 (.D(mem_rdata_7__N_185[20]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i20.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i19 (.D(mem_rdata_7__N_185[19]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i19.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i18 (.D(mem_rdata_7__N_185[18]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i18.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i13 (.D(mem_rdata_7__N_185[13]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i13.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i12 (.D(mem_rdata_7__N_185[12]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i12.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i11 (.D(mem_rdata_7__N_185[11]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i11.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i10 (.D(mem_rdata_7__N_185[10]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i10.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i9 (.D(mem_rdata_7__N_185[9]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i9.GSR = "DISABLED";
    FD1P3IX spi_sdo_r__i8 (.D(mem_rdata_7__N_185[8]), .SP(clk_enable_523), 
            .CD(n29239), .CK(clk), .Q(spi_sdo_r[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i8.GSR = "DISABLED";
    FD1P3AX spi_sdo_r__i7 (.D(n27172), .SP(clk_enable_523), .CK(clk), 
            .Q(spi_sdo_r[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i7.GSR = "DISABLED";
    FD1P3AX spi_sdo_r__i6 (.D(n27179), .SP(clk_enable_523), .CK(clk), 
            .Q(spi_sdo_r[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i6.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(n35), .B(spi_sdo_valid_N_297), .C(n40), .D(n36), 
         .Z(spi_sdo_39__N_145[2])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(\spi_data_out_r_39__N_2643[2] ), .B(n28), .C(n13), 
         .D(clear_intrpt), .Z(n35)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i14_4_lut.init = 16'hfefc;
    LUT4 i19_4_lut (.A(n31_c), .B(n38), .C(n4), .D(n22), .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i15_4_lut (.A(\spi_data_out_r_39__N_934[2] ), .B(n30), .C(n19), 
         .D(spi_data_out_r_39__N_974), .Z(n36)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i15_4_lut.init = 16'hfefc;
    FD1P3IX spi_data_valid_r_58 (.D(spi_data_valid), .SP(clk_enable_341), 
            .CD(n29247), .CK(clk), .Q(spi_data_valid_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_valid_r_58.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i1 (.D(spi_cmd[1]), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(spi_cmd_r[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i1.GSR = "DISABLED";
    LUT4 i7_4_lut (.A(\spi_data_out_r_39__N_4157[2] ), .B(\spi_data_out_r_39__N_1168[2] ), 
         .C(spi_data_out_r_39__N_4197), .D(spi_data_out_r_39__N_1208), .Z(n28)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i7_4_lut.init = 16'heca0;
    LUT4 i10_4_lut (.A(\spi_data_out_r_39__N_2927[2] ), .B(\spi_data_out_r_39__N_2785[2] ), 
         .C(clear_intrpt_adj_151), .D(clear_intrpt_adj_152), .Z(n31_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i10_4_lut.init = 16'heca0;
    LUT4 i17_4_lut (.A(n8), .B(n34), .C(n24_c), .D(n15), .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i17_4_lut.init = 16'hfffe;
    FD1P3IX spi_cmd_r__i2 (.D(spi_cmd[2]), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(spi_cmd_r[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i2.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i3 (.D(spi_cmd_c[3]), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(spi_cmd_r[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i3.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i4 (.D(\spi_cmd[4] ), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(spi_cmd_r_c[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i4.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i5 (.D(spi_cmd_c[5]), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(spi_cmd_r_c[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i5.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i6 (.D(spi_cmd_c[6]), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(\spi_cmd_r[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i6.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i7 (.D(spi_cmd_c[7]), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(\spi_cmd_r[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i7.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i8 (.D(spi_cmd_c[8]), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(\spi_cmd_r[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i8.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i9 (.D(spi_cmd_c[9]), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(\spi_cmd_r[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i9.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i10 (.D(spi_cmd_c[10]), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(\spi_cmd_r[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i10.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i11 (.D(spi_cmd_c[11]), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(\spi_cmd_r[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i11.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i12 (.D(spi_cmd_c[12]), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(\spi_cmd_r[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i12.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i13 (.D(spi_cmd_c[13]), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(\spi_cmd_r[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i13.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i14 (.D(spi_cmd_c[14]), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(\spi_cmd_r[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i14.GSR = "DISABLED";
    FD1P3IX spi_cmd_r__i15 (.D(\spi_cmd[15] ), .SP(clk_enable_357), .CD(n29247), 
            .CK(clk), .Q(\spi_cmd_r[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_cmd_r__i15.GSR = "DISABLED";
    FD1P3AX spi_sdo_r__i5 (.D(n27173), .SP(clk_enable_523), .CK(clk), 
            .Q(spi_sdo_r[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i5.GSR = "DISABLED";
    FD1P3IX spi_sdo__i1 (.D(\spi_data_out_r[1] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i1.GSR = "DISABLED";
    FD1P3IX spi_sdo__i3 (.D(\spi_data_out_r[3] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i3.GSR = "DISABLED";
    FD1P3IX spi_sdo__i4 (.D(\spi_data_out_r[4] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i4.GSR = "DISABLED";
    FD1P3IX spi_sdo__i5 (.D(\spi_data_out_r[5] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i5.GSR = "DISABLED";
    FD1P3IX spi_sdo__i6 (.D(\spi_data_out_r[6] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i6.GSR = "DISABLED";
    FD1P3IX spi_sdo__i7 (.D(\spi_data_out_r[7] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i7.GSR = "DISABLED";
    FD1P3IX spi_sdo__i8 (.D(\spi_data_out_r[8] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i8.GSR = "DISABLED";
    FD1P3IX spi_sdo__i9 (.D(\spi_data_out_r[9] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i9.GSR = "DISABLED";
    FD1P3IX spi_sdo__i10 (.D(\spi_data_out_r[10] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i10.GSR = "DISABLED";
    FD1P3IX spi_sdo__i11 (.D(\spi_data_out_r[11] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i11.GSR = "DISABLED";
    FD1P3IX spi_sdo__i12 (.D(\spi_data_out_r[12] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i12.GSR = "DISABLED";
    FD1P3IX spi_sdo__i13 (.D(\spi_data_out_r[13] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i13.GSR = "DISABLED";
    FD1P3IX spi_sdo__i14 (.D(\spi_data_out_r[14] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i14.GSR = "DISABLED";
    FD1P3IX spi_sdo__i15 (.D(\spi_data_out_r[15] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i15.GSR = "DISABLED";
    FD1P3IX spi_sdo__i16 (.D(\spi_data_out_r[16] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i16.GSR = "DISABLED";
    FD1P3IX spi_sdo__i17 (.D(\spi_data_out_r[17] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i17.GSR = "DISABLED";
    FD1P3IX spi_sdo__i18 (.D(\spi_data_out_r[18] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i18.GSR = "DISABLED";
    FD1P3IX spi_sdo__i19 (.D(\spi_data_out_r[19] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i19.GSR = "DISABLED";
    FD1P3IX spi_sdo__i20 (.D(\spi_data_out_r[20] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i20.GSR = "DISABLED";
    FD1P3IX spi_sdo__i21 (.D(\spi_data_out_r[21] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i21.GSR = "DISABLED";
    FD1P3IX spi_sdo__i22 (.D(\spi_data_out_r[22] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i22.GSR = "DISABLED";
    FD1P3IX spi_sdo__i23 (.D(\spi_data_out_r[23] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i23.GSR = "DISABLED";
    FD1P3IX spi_sdo__i24 (.D(\spi_data_out_r[24] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i24.GSR = "DISABLED";
    FD1P3IX spi_sdo__i25 (.D(\spi_data_out_r[25] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i25.GSR = "DISABLED";
    FD1P3IX spi_sdo__i26 (.D(\spi_data_out_r[26] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i26.GSR = "DISABLED";
    FD1P3IX spi_sdo__i27 (.D(\spi_data_out_r[27] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i27.GSR = "DISABLED";
    FD1P3IX spi_sdo__i28 (.D(\spi_data_out_r[28] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i28.GSR = "DISABLED";
    FD1P3IX spi_sdo__i29 (.D(\spi_data_out_r[29] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i29.GSR = "DISABLED";
    FD1P3IX spi_sdo__i30 (.D(\spi_data_out_r[30] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i30.GSR = "DISABLED";
    FD1P3IX spi_sdo__i31 (.D(\spi_data_out_r[31] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i31.GSR = "DISABLED";
    FD1P3IX spi_sdo__i32 (.D(\spi_data_out_r[32] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i32.GSR = "DISABLED";
    FD1P3IX spi_sdo__i33 (.D(\spi_data_out_r[33] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i33.GSR = "DISABLED";
    FD1P3IX spi_sdo__i34 (.D(\spi_data_out_r[34] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i34.GSR = "DISABLED";
    FD1P3IX spi_sdo__i35 (.D(\spi_data_out_r[35] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i35.GSR = "DISABLED";
    FD1P3IX spi_sdo__i36 (.D(\spi_data_out_r[36] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i36.GSR = "DISABLED";
    FD1P3IX spi_sdo__i37 (.D(\spi_data_out_r[37] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i37.GSR = "DISABLED";
    FD1P3IX spi_sdo__i38 (.D(\spi_data_out_r[38] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i38.GSR = "DISABLED";
    FD1P3IX spi_sdo__i39 (.D(\spi_data_out_r[39] ), .SP(spi_sdo_valid_N_296), 
            .CD(n10988), .CK(clk), .Q(spi_sdo[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(91[9] 108[5])
    defparam spi_sdo__i39.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_566 (.A(\spi_data_out_r_39__N_5174[2] ), .B(\spi_data_out_r_39__N_3818[2] ), 
         .C(spi_data_out_r_39__N_5214), .D(spi_data_out_r_39__N_3858), .Z(n22)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i1_4_lut_adj_566.init = 16'heca0;
    LUT4 i13_4_lut (.A(\spi_data_out_r_39__N_5852[2] ), .B(n26_c), .C(n11), 
         .D(spi_data_out_r_39__N_5892), .Z(n34)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i13_4_lut.init = 16'hfefc;
    LUT4 i3_4_lut_adj_567 (.A(\spi_data_out_r_39__N_4496[2] ), .B(\spi_data_out_r_39__N_1870[2] ), 
         .C(spi_data_out_r_39__N_4536), .D(spi_data_out_r_39__N_1910), .Z(n24_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i3_4_lut_adj_567.init = 16'heca0;
    LUT4 i5_4_lut (.A(\spi_data_out_r_39__N_5513[2] ), .B(\spi_data_out_r_39__N_1636[2] ), 
         .C(spi_data_out_r_39__N_5553), .D(spi_data_out_r_39__N_1676), .Z(n26_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i5_4_lut.init = 16'heca0;
    LUT4 i9_4_lut (.A(\spi_data_out_r_39__N_2104[2] ), .B(\spi_data_out_r_39__N_2572[2] ), 
         .C(spi_data_out_r_39__N_2144), .D(clear_intrpt_adj_153), .Z(n30)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i9_4_lut.init = 16'heca0;
    LUT4 i1_2_lut_rep_583 (.A(spi_cmd_r_c[5]), .B(spi_cmd_r_c[4]), .Z(n29311)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_583.init = 16'h8888;
    LUT4 i1_2_lut_rep_446_3_lut (.A(spi_cmd_r_c[5]), .B(spi_cmd_r_c[4]), 
         .C(spi_cmd_r[0]), .Z(n29174)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_446_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_488_3_lut (.A(spi_cmd_r_c[5]), .B(spi_cmd_r_c[4]), 
         .C(spi_cmd_r[3]), .Z(n29216)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_488_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_rep_346_3_lut_4_lut (.A(\spi_addr_r[1] ), .B(n29121), 
         .C(spi_cmd_r[2]), .D(n29182), .Z(n29074)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_346_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_347_3_lut_4_lut (.A(\spi_addr_r[1] ), .B(n29121), 
         .C(n27058), .D(n29182), .Z(n29075)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_347_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_350_3_lut_4_lut (.A(\spi_addr_r[1] ), .B(n29121), 
         .C(n29174), .D(spi_cmd_r[2]), .Z(n29078)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_350_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_351_3_lut_4_lut (.A(\spi_addr_r[1] ), .B(n29121), 
         .C(n27259), .D(spi_cmd_r[2]), .Z(n29079)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_351_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_352_3_lut_4_lut (.A(\spi_addr_r[1] ), .B(n29121), 
         .C(n29162), .D(spi_cmd_r[2]), .Z(n29080)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_352_3_lut_4_lut.init = 16'h0040;
    LUT4 mux_18_i15_3_lut (.A(spi_sdo_r[6]), .B(spi_sdo[14]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i15_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_344_3_lut_4_lut (.A(spi_cmd_r[2]), .B(n29121), .C(n29254), 
         .D(n27286), .Z(n29072)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_344_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_rep_343_3_lut_4_lut (.A(spi_cmd_r[2]), .B(n29121), .C(n65_adj_154), 
         .D(n27286), .Z(n29071)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_343_3_lut_4_lut.init = 16'h4000;
    LUT4 i2_3_lut_rep_364_4_lut (.A(spi_cmd_r[2]), .B(n29121), .C(n29162), 
         .D(\spi_addr_r[1] ), .Z(n29092)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i2_3_lut_rep_364_4_lut.init = 16'h4000;
    LUT4 i1_4_lut_adj_568 (.A(n37), .B(spi_sdo_valid_N_297), .C(n42), 
         .D(n38_adj_6731), .Z(spi_sdo_39__N_145[0])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i1_4_lut_adj_568.init = 16'hfffe;
    LUT4 i15_4_lut_adj_569 (.A(\spi_data_out_r_39__N_2927[0] ), .B(n30_adj_6732), 
         .C(n17), .D(clear_intrpt_adj_151), .Z(n37)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i15_4_lut_adj_569.init = 16'hfefc;
    LUT4 i20_4_lut (.A(n3), .B(n40_adj_6733), .C(n34_adj_6734), .D(n20), 
         .Z(n42)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i16_4_lut (.A(\spi_data_out_r_39__N_3818[0] ), .B(n32_c), .C(n4_adj_155), 
         .D(spi_data_out_r_39__N_3858), .Z(n38_adj_6731)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i16_4_lut.init = 16'hfefc;
    LUT4 i8_4_lut (.A(\spi_data_out_r_39__N_1870[0] ), .B(\spi_data_out_r_39__N_2785[0] ), 
         .C(spi_data_out_r_39__N_1910), .D(clear_intrpt_adj_152), .Z(n30_adj_6732)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i8_4_lut.init = 16'heca0;
    LUT4 i18_4_lut (.A(n15_adj_156), .B(n36_adj_6737), .C(n26_adj_6738), 
         .D(n2), .Z(n40_adj_6733)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i12_4_lut (.A(\spi_data_out_r_39__N_4496[0] ), .B(n24_adj_6739), 
         .C(n11_adj_157), .D(spi_data_out_r_39__N_4536), .Z(n34_adj_6734)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i12_4_lut.init = 16'hfefc;
    LUT4 i14_4_lut_adj_570 (.A(\spi_data_out_r_39__N_4835[0] ), .B(n28_adj_6741), 
         .C(n21), .D(spi_data_out_r_39__N_4875), .Z(n36_adj_6737)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i14_4_lut_adj_570.init = 16'hfefc;
    LUT4 i4_4_lut (.A(\spi_data_out_r_39__N_770[0] ), .B(\spi_data_out_r_39__N_5852[0] ), 
         .C(spi_data_out_r_39__N_810), .D(spi_data_out_r_39__N_5892), .Z(n26_adj_6738)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i4_4_lut.init = 16'heca0;
    LUT4 i6_4_lut (.A(\spi_data_out_r_39__N_2338[0] ), .B(\spi_data_out_r_39__N_2572[0] ), 
         .C(spi_data_out_r_39__N_2378), .D(clear_intrpt_adj_153), .Z(n28_adj_6741)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i6_4_lut.init = 16'heca0;
    LUT4 i10_4_lut_adj_571 (.A(\spi_data_out_r_39__N_2104[0] ), .B(\spi_data_out_r_39__N_2856[0] ), 
         .C(spi_data_out_r_39__N_2144), .D(clear_intrpt_adj_158), .Z(n32_c)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i10_4_lut_adj_571.init = 16'heca0;
    LUT4 i2_4_lut (.A(\spi_data_out_r_39__N_1636[0] ), .B(\spi_data_out_r_39__N_2643[0] ), 
         .C(spi_data_out_r_39__N_1676), .D(clear_intrpt), .Z(n24_adj_6739)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_slave_top.v(100[8] 107[6])
    defparam i2_4_lut.init = 16'heca0;
    LUT4 mux_18_i40_3_lut (.A(spi_sdo_r[31]), .B(spi_sdo[39]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[39])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i40_3_lut.init = 16'hcaca;
    LUT4 mux_18_i39_3_lut (.A(spi_sdo_r[30]), .B(spi_sdo[38]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[38])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i39_3_lut.init = 16'hcaca;
    LUT4 mux_18_i38_3_lut (.A(spi_sdo_r[29]), .B(spi_sdo[37]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[37])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i38_3_lut.init = 16'hcaca;
    LUT4 mux_18_i37_3_lut (.A(spi_sdo_r[28]), .B(spi_sdo[36]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[36])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i37_3_lut.init = 16'hcaca;
    LUT4 mux_18_i36_3_lut (.A(spi_sdo_r[27]), .B(spi_sdo[35]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[35])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i36_3_lut.init = 16'hcaca;
    LUT4 mux_18_i35_3_lut (.A(spi_sdo_r[26]), .B(spi_sdo[34]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[34])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i35_3_lut.init = 16'hcaca;
    LUT4 mux_18_i34_3_lut (.A(spi_sdo_r[25]), .B(spi_sdo[33]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[33])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i34_3_lut.init = 16'hcaca;
    LUT4 mux_18_i33_3_lut (.A(spi_sdo_r[24]), .B(spi_sdo[32]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[32])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i33_3_lut.init = 16'hcaca;
    LUT4 mux_18_i32_3_lut (.A(spi_sdo_r[23]), .B(spi_sdo[31]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i32_3_lut.init = 16'hcaca;
    LUT4 mux_18_i31_3_lut (.A(spi_sdo_r[22]), .B(spi_sdo[30]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i31_3_lut.init = 16'hcaca;
    LUT4 mux_18_i30_3_lut (.A(spi_sdo_r[21]), .B(spi_sdo[29]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i30_3_lut.init = 16'hcaca;
    LUT4 mux_18_i29_3_lut (.A(spi_sdo_r[20]), .B(spi_sdo[28]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i29_3_lut.init = 16'hcaca;
    LUT4 mux_18_i28_3_lut (.A(spi_sdo_r[19]), .B(spi_sdo[27]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i28_3_lut.init = 16'hcaca;
    LUT4 mux_18_i27_3_lut (.A(spi_sdo_r[18]), .B(spi_sdo[26]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i27_3_lut.init = 16'hcaca;
    LUT4 mux_18_i26_3_lut (.A(spi_sdo_r[17]), .B(spi_sdo[25]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i26_3_lut.init = 16'hcaca;
    LUT4 mux_18_i25_3_lut (.A(spi_sdo_r[16]), .B(spi_sdo[24]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i25_3_lut.init = 16'hcaca;
    LUT4 mux_18_i24_3_lut (.A(spi_sdo_r[15]), .B(spi_sdo[23]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i24_3_lut.init = 16'hcaca;
    LUT4 mux_18_i23_3_lut (.A(spi_sdo_r[14]), .B(spi_sdo[22]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i23_3_lut.init = 16'hcaca;
    LUT4 mux_18_i22_3_lut (.A(spi_sdo_r[13]), .B(spi_sdo[21]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i22_3_lut.init = 16'hcaca;
    LUT4 mux_18_i21_3_lut (.A(spi_sdo_r[12]), .B(spi_sdo[20]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i21_3_lut.init = 16'hcaca;
    LUT4 mux_18_i20_3_lut (.A(spi_sdo_r[11]), .B(spi_sdo[19]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i20_3_lut.init = 16'hcaca;
    LUT4 mux_18_i19_3_lut (.A(spi_sdo_r[10]), .B(spi_sdo[18]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i19_3_lut.init = 16'hcaca;
    LUT4 mux_18_i14_3_lut (.A(spi_sdo_r[5]), .B(spi_sdo[13]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i14_3_lut.init = 16'hcaca;
    LUT4 mux_18_i13_3_lut (.A(spi_sdo_r[4]), .B(spi_sdo[12]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i13_3_lut.init = 16'hcaca;
    LUT4 mux_18_i12_3_lut (.A(spi_sdo_r[3]), .B(spi_sdo[11]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i12_3_lut.init = 16'hcaca;
    LUT4 mux_18_i11_3_lut (.A(spi_sdo_r[2]), .B(spi_sdo[10]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i11_3_lut.init = 16'hcaca;
    LUT4 mux_18_i10_3_lut (.A(spi_sdo_r[1]), .B(spi_sdo[9]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i10_3_lut.init = 16'hcaca;
    LUT4 mux_18_i9_3_lut (.A(spi_sdo_r[0]), .B(spi_sdo[8]), .C(spi_sdo_valid), 
         .Z(mem_rdata_7__N_185[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_slave_top.v(116[8] 119[27])
    defparam mux_18_i9_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_572 (.A(\spi_addr_r[2] ), .B(spi_cmd_r[2]), .Z(n60)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_adj_572.init = 16'h4444;
    LUT4 i1_3_lut_4_lut (.A(n29089), .B(n65_adj_154), .C(n27338), .D(n13074), 
         .Z(clk_enable_206)) /* synthesis lut_function=(A (B (C+!(D)))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_3_lut_4_lut.init = 16'h8088;
    LUT4 i1_2_lut_rep_358_3_lut_4_lut (.A(n29130), .B(\spi_addr_r[2] ), 
         .C(n29182), .D(\spi_addr_r[1] ), .Z(n29086)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_358_3_lut_4_lut.init = 16'h0008;
    LUT4 spi_addr_valid_r_I_5_3_lut (.A(spi_sdo_valid_N_296), .B(spi_addr_valid), 
         .C(spi_data_valid), .Z(spi_addr_valid_r_N_303)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // c:/s_links/sources/mcm_top.v(186[3] 206[2])
    defparam spi_addr_valid_r_I_5_3_lut.init = 16'hecec;
    LUT4 i1_2_lut_rep_362_3_lut_4_lut (.A(n29130), .B(\spi_addr_r[2] ), 
         .C(spi_cmd_r[2]), .D(\spi_addr_r[1] ), .Z(n29090)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_362_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_rep_361_3_lut_4_lut (.A(n29130), .B(\spi_addr_r[2] ), 
         .C(n27286), .D(spi_cmd_r[2]), .Z(n29089)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_361_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_368_3_lut_4_lut (.A(n29169), .B(n29182), .C(resetn_c), 
         .D(n29127), .Z(n29096)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_368_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_369_3_lut_4_lut (.A(n29169), .B(n29182), .C(n29213), 
         .D(n29127), .Z(n29097)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_369_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_378_3_lut_4_lut (.A(n29169), .B(n29182), .C(n13074), 
         .D(n29127), .Z(n29106)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_378_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_379_3_lut_4_lut (.A(n27), .B(n29144), .C(\spi_addr_r[1] ), 
         .D(\spi_addr_r[2] ), .Z(n29107)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_379_3_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_rep_383_3_lut_4_lut (.A(n27), .B(n29144), .C(spi_cmd_r[2]), 
         .D(\spi_addr_r[2] ), .Z(n29111)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i1_2_lut_rep_383_3_lut_4_lut.init = 16'h0400;
    LUT4 i2_3_lut_rep_395_4_lut (.A(n27), .B(n29144), .C(n29251), .D(spi_cmd_r[0]), 
         .Z(n29123)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam i2_3_lut_rep_395_4_lut.init = 16'h0004;
    FD1P3AX spi_sdo_r__i4 (.D(n27174), .SP(clk_enable_523), .CK(clk), 
            .Q(spi_sdo_r[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i4.GSR = "DISABLED";
    FD1P3AX spi_sdo_r__i3 (.D(n27175), .SP(clk_enable_523), .CK(clk), 
            .Q(spi_sdo_r[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(111[11] 120[7])
    defparam spi_sdo_r__i3.GSR = "DISABLED";
    FD1P3IX spi_data_r__i0_rep_594 (.D(spi_data[0]), .SP(clk_enable_524), 
            .CD(n29247), .CK(clk), .Q(n29762)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=186, LSE_RLINE=206 */ ;   // c:/s_links/sources/spi_slave_top.v(123[11] 150[5])
    defparam spi_data_r__i0_rep_594.GSR = "DISABLED";
    wb_ctrl wb_ctrl_inst (.wb_cyc_i(wb_cyc_i), .clk(clk), .clk_enable_95(clk_enable_95), 
            .wb_cyc_i_N_339(wb_cyc_i_N_339), .\wb_adr_i[0] (wb_adr_i[0]), 
            .\address[0] (address[0]), .wb_we_i(wb_we_i), .wb_we_i_N_344(wb_we_i_N_344), 
            .wb_dat_i({wb_dat_i}), .wr_data({wr_data}), .wb_sm(wb_sm), 
            .n28767(n28767), .n29268(n29268), .\address_7__N_549[1] (address_7__N_549[1]), 
            .spi_cmd_start(spi_cmd_start), .\address_7__N_565[1] (address_7__N_565[1]), 
            .\wb_adr_i[1] (wb_adr_i[1]), .\address[1] (address[1]), .\wb_adr_i[4] (wb_adr_i[4]), 
            .n29757(n29757), .wr_en(wr_en), .wr_en_N_355(wr_en_N_355)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/spi_slave_top.v(179[12] 196[15])
    spi_slave_efb spi_slave_efb_inst (.clk(clk), .n29239(n29239), .wb_cyc_i(wb_cyc_i), 
            .wb_we_i(wb_we_i), .GND_net(GND_net), .\wb_adr_i[4] (wb_adr_i[4]), 
            .\wb_adr_i[1] (wb_adr_i[1]), .\wb_adr_i[0] (wb_adr_i[0]), .wb_dat_i({wb_dat_i}), 
            .spi_scsn_c(spi_scsn_c), .wb_dat_o({wb_dat_o}), .\address_7__N_549[1] (address_7__N_549[1]), 
            .spi_mosi_oe(spi_mosi_oe), .spi_mosi_o(spi_mosi_o), .spi_miso_oe(spi_miso_oe), 
            .spi_miso_o(spi_miso_o), .spi_clk_oe(spi_clk_oe), .spi_clk_o(spi_clk_o), 
            .spi_mosi_i(spi_mosi_i), .spi_miso_i(spi_miso_i), .spi_clk_i(spi_clk_i), 
            .VCC_net(VCC_net), .n2720(n2713[9]), .mem_rdata_update_N_729(mem_rdata_update_N_729), 
            .spi_addr_valid_N_732(spi_addr_valid_N_732), .n29176(n29176), 
            .n2724(n2713[5]), .n29179(n29179), .n7083(n7083), .clk_enable_309(clk_enable_309), 
            .clk_enable_516(clk_enable_516), .wb_sm(wb_sm), .clk_enable_95(clk_enable_95)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/s_links/sources/spi_slave_top.v(162[18] 176[15])
    spi_ctrl spi_ctrl_inst (.spi_addr_valid(spi_addr_valid), .clk(clk), 
            .spi_addr_valid_N_732(spi_addr_valid_N_732), .clk_enable_516(clk_enable_516), 
            .n29176(n29176), .\address_7__N_549[1] (address_7__N_549[1]), 
            .mem_rdata_update_N_729(mem_rdata_update_N_729), .resetn_c(resetn_c), 
            .n29239(n29239), .quad_set_complete(quad_set_complete), .n29162(n29162), 
            .n29090(n29090), .clk_enable_518(clk_enable_518), .spi_sdo_valid(spi_sdo_valid), 
            .clk_enable_523(clk_enable_523), .n29127(n29127), .n29211(n29211), 
            .n27225(n27225), .clk_enable_398(clk_enable_398), .n29254(n29254), 
            .n29102(n29102), .n29255(n29255), .clk_enable_188(clk_enable_188), 
            .n6(n6), .clk_enable_303(clk_enable_303), .n32(n32), .\quad_homing[1] (\quad_homing[1] ), 
            .n27657(n27657), .n24(n24), .n27201(n27201), .n60(n60), 
            .n29123(n29123), .clk_enable_179(clk_enable_179), .n29213(n29213), 
            .\spi_cmd_r[2] (spi_cmd_r[2]), .n29086(n29086), .clk_enable_182(clk_enable_182), 
            .clear_intrpt(clear_intrpt_adj_152), .intrpt_out_N_2848(intrpt_out_N_2848), 
            .n29100(n29100), .clk_enable_185(clk_enable_185), .wr_data({wr_data}), 
            .n29134(n29134), .n27280(n27280), .clk_enable_509(clk_enable_509), 
            .reset_r_N_4813(reset_r_N_4813), .EM_STOP(EM_STOP), .n29070(n29070), 
            .clk_enable_306(clk_enable_306), .n29101(n29101), .\spi_addr_r[2] (\spi_addr_r[2] ), 
            .clk_enable_186(clk_enable_186), .quad_set_complete_adj_135(quad_set_complete_adj_159), 
            .n29120(n29120), .clk_enable_505(clk_enable_505), .\spi_addr_r[1] (\spi_addr_r[1] ), 
            .n29111(n29111), .clk_enable_76(clk_enable_76), .n29104(n29104), 
            .\spi_cmd_r[3] (spi_cmd_r[3]), .clk_enable_436(clk_enable_436), 
            .n19233(n19233), .clk_enable_184(clk_enable_184), .n29129(n29129), 
            .clk_enable_204(clk_enable_204), .clear_intrpt_adj_136(clear_intrpt_adj_153), 
            .intrpt_out_N_2635(intrpt_out_N_2635), .n29288(n29288), .clk_enable_183(clk_enable_183), 
            .n29095(n29095), .clk_enable_271(clk_enable_271), .n29072(n29072), 
            .n29083(n29083), .clk_enable_521(clk_enable_521), .quad_set_valid(quad_set_valid), 
            .n66(n66), .n21446(n21446), .clk_1MHz_enable_171(clk_1MHz_enable_171), 
            .n29124(n29124), .clk_enable_197(clk_enable_197), .n26948(n26948), 
            .n13(n13_adj_160), .n12714(n12714), .n27301(n27301), .n29242(n29242), 
            .clk_enable_193(clk_enable_193), .\spi_cmd_r[0] (spi_cmd_r[0]), 
            .n29074(n29074), .clk_enable_200(clk_enable_200), .spi_sdo_valid_N_297(spi_sdo_valid_N_297), 
            .n10988(n10988), .n29307(n29307), .n27286(n27286), .clk_enable_499(clk_enable_499), 
            .n4(n4_c), .n27240(n27240), .clk_enable_32(clk_enable_32), 
            .quad_set_complete_adj_137(quad_set_complete_adj_161), .n29092(n29092), 
            .clk_enable_520(clk_enable_520), .n29286(n29286), .clk_enable_77(clk_enable_77), 
            .clear_intrpt_adj_138(clear_intrpt), .intrpt_out_N_2706(intrpt_out_N_2706), 
            .quad_set_valid_adj_139(quad_set_valid_adj_162), .n79(n79), 
            .n20819(n20819), .clk_1MHz_enable_340(clk_1MHz_enable_340), 
            .n27285(n27285), .n29110(n29110), .clk_enable_340(clk_enable_340), 
            .n31(n31), .\quad_homing[1]_adj_140 (\quad_homing[1]_adj_163 ), 
            .n5(n5), .n26(n26), .n27234(n27234), .clk_enable_174(clk_enable_174), 
            .n27243(n27243), .clk_enable_171(clk_enable_171), .clk_enable_172(clk_enable_172), 
            .n29119(n29119), .n29174(n29174), .clk_enable_435(clk_enable_435), 
            .n29082(n29082), .n29106(n29106), .clk_enable_506(clk_enable_506), 
            .\spi_data[0] (spi_data[0]), .wb_dat_o({wb_dat_o}), .n29144(n29144), 
            .clk_enable_269(clk_enable_269), .n13074(n13074), .clk_enable_167(clk_enable_167), 
            .n29175(n29175), .clk_enable_28(clk_enable_28), .clk_enable_309(clk_enable_309), 
            .n29179(n29179), .n27259(n27259), .n29107(n29107), .clk_enable_131(clk_enable_131), 
            .clear_intrpt_adj_141(clear_intrpt_adj_158), .intrpt_out_N_2919(intrpt_out_N_2919), 
            .n65(n65), .clk_enable_194(clk_enable_194), .n65_adj_142(n65_adj_154), 
            .clk_enable_177(clk_enable_177), .spi_sdo_valid_N_296(spi_sdo_valid_N_296), 
            .clk_enable_305(clk_enable_305), .clk_enable_189(clk_enable_189), 
            .\address[0] (address[0]), .clk_enable_180(clk_enable_180), 
            .wr_en(wr_en), .spi_scsn_c(spi_scsn_c), .clk_enable_162(clk_enable_162), 
            .clk_enable_166(clk_enable_166), .n29256(n29256), .clk_enable_175(clk_enable_175), 
            .clk_enable_176(clk_enable_176), .quad_set_complete_adj_143(quad_set_complete_adj_164), 
            .n29105(n29105), .clk_enable_502(clk_enable_502), .n29071(n29071), 
            .n29077(n29077), .clk_enable_526(clk_enable_526), .n29069(n29069), 
            .n29075(n29075), .clk_enable_342(clk_enable_342), .clk_enable_202(clk_enable_202), 
            .clear_intrpt_adj_144(clear_intrpt_adj_151), .intrpt_out_N_2990(intrpt_out_N_2990), 
            .clk_enable_201(clk_enable_201), .clk_enable_467(clk_enable_467), 
            .clk_enable_191(clk_enable_191), .clk_enable_187(clk_enable_187), 
            .clk_enable_192(clk_enable_192), .quad_set_complete_adj_145(quad_set_complete_adj_165), 
            .clk_enable_519(clk_enable_519), .clk_enable_170(clk_enable_170), 
            .n29118(n29118), .n29214(n29214), .clk_enable_286(clk_enable_286), 
            .n29182(n29182), .clk_enable_359(clk_enable_359), .reset_r_N_4474(reset_r_N_4474), 
            .n29097(n29097), .clk_enable_307(clk_enable_307), .clear_intrpt_adj_146(clear_intrpt_adj_166), 
            .intrpt_out_N_3061(intrpt_out_N_3061), .clk_enable_86(clk_enable_86), 
            .clk_enable_181(clk_enable_181), .clk_enable_288(clk_enable_288), 
            .clk_enable_433(clk_enable_433), .clk_enable_434(clk_enable_434), 
            .quad_set_complete_adj_147(quad_set_complete_adj_167), .clk_enable_501(clk_enable_501), 
            .n29205(n29205), .clk_enable_169(clk_enable_169), .clear_intrpt_adj_148(clear_intrpt_adj_168), 
            .intrpt_out_N_2777(intrpt_out_N_2777), .n27058(n27058), .clk_enable_400(clk_enable_400), 
            .clk_enable_402(clk_enable_402), .quad_set_complete_adj_149(quad_set_complete_adj_169), 
            .clk_enable_503(clk_enable_503), .clk_enable_30(clk_enable_30), 
            .n2724(n2713[5]), .n2720(n2713[9]), .spi_cmd({\spi_cmd[15] , 
            spi_cmd_c[14:5], \spi_cmd[4] , spi_cmd_c[3], spi_cmd[2:1], 
            \spi_cmd[0] }), .wr_en_N_355(wr_en_N_355), .n9633(n9633), 
            .spi_addr({spi_addr_c[7:4], \spi_addr[3] , \spi_addr[2] , 
            \spi_addr[1] , spi_addr[0]}), .n27465(n27465), .n26928(n26928), 
            .n29141(n29141), .n29126(n29126), .n27618(n27618), .spi_cmd_start(spi_cmd_start), 
            .n29268(n29268), .wb_sm(wb_sm), .n28767(n28767), .wb_cyc_i_N_339(wb_cyc_i_N_339), 
            .\address_7__N_565[1] (address_7__N_565[1]), .n7083(n7083), 
            .mem_rdata({mem_rdata}), .GND_net(GND_net), .n29114(n29114), 
            .clk_enable_20(clk_enable_20), .\spi_data[1] (spi_data[1]), 
            .\spi_data[2] (spi_data[2]), .\spi_data[3] (spi_data[3]), .\spi_data[4] (spi_data[4]), 
            .\spi_data[5] (spi_data[5]), .\spi_data[6] (spi_data[6]), .\spi_data[7] (spi_data[7]), 
            .\spi_data[8] (spi_data[8]), .\spi_data[9] (spi_data[9]), .\spi_data[10] (spi_data[10]), 
            .\spi_data[11] (spi_data[11]), .\spi_data[12] (spi_data[12]), 
            .\spi_data[13] (spi_data[13]), .\spi_data[14] (spi_data[14]), 
            .\spi_data[15] (spi_data[15]), .\spi_data[16] (spi_data[16]), 
            .\spi_data[17] (spi_data[17]), .\spi_data[18] (spi_data[18]), 
            .\spi_data[19] (spi_data[19]), .\spi_data[20] (spi_data[20]), 
            .\spi_data[21] (spi_data[21]), .\spi_data[22] (spi_data[22]), 
            .\spi_data[23] (spi_data[23]), .\spi_data[24] (spi_data[24]), 
            .\spi_data[25] (spi_data[25]), .\spi_data[26] (spi_data[26]), 
            .\spi_data[27] (spi_data[27]), .\spi_data[28] (spi_data[28]), 
            .\spi_data[29] (spi_data[29]), .\spi_data[30] (spi_data[30]), 
            .\spi_data[31] (spi_data[31]), .\address[1] (address[1]), .spi_data_valid(spi_data_valid), 
            .spi_cmd_valid(spi_cmd_valid), .n31_adj_150(n31_adj_170), .wb_we_i_N_344(wb_we_i_N_344), 
            .n29761(n29761)) /* synthesis syn_module_defined=1 */ ;   // c:/s_links/sources/spi_slave_top.v(203[4] 225[21])
    
endmodule
//
// Verilog Description of module wb_ctrl
//

module wb_ctrl (wb_cyc_i, clk, clk_enable_95, wb_cyc_i_N_339, \wb_adr_i[0] , 
            \address[0] , wb_we_i, wb_we_i_N_344, wb_dat_i, wr_data, 
            wb_sm, n28767, n29268, \address_7__N_549[1] , spi_cmd_start, 
            \address_7__N_565[1] , \wb_adr_i[1] , \address[1] , \wb_adr_i[4] , 
            n29757, wr_en, wr_en_N_355) /* synthesis syn_module_defined=1 */ ;
    output wb_cyc_i;
    input clk;
    input clk_enable_95;
    input wb_cyc_i_N_339;
    output \wb_adr_i[0] ;
    input \address[0] ;
    output wb_we_i;
    input wb_we_i_N_344;
    output [7:0]wb_dat_i;
    input [7:0]wr_data;
    output wb_sm;
    input n28767;
    input n29268;
    input \address_7__N_549[1] ;
    input spi_cmd_start;
    output \address_7__N_565[1] ;
    output \wb_adr_i[1] ;
    input \address[1] ;
    output \wb_adr_i[4] ;
    input n29757;
    input wr_en;
    output wr_en_N_355;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    FD1P3AX wb_cyc_i_36 (.D(wb_cyc_i_N_339), .SP(clk_enable_95), .CK(clk), 
            .Q(wb_cyc_i)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_cyc_i_36.GSR = "ENABLED";
    FD1P3AX wb_adr_i_i0 (.D(\address[0] ), .SP(wb_cyc_i_N_339), .CK(clk), 
            .Q(\wb_adr_i[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_adr_i_i0.GSR = "ENABLED";
    FD1P3AX wb_we_i_38 (.D(wb_we_i_N_344), .SP(clk_enable_95), .CK(clk), 
            .Q(wb_we_i)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_we_i_38.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i0 (.D(wr_data[0]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i0.GSR = "ENABLED";
    FD1S3AX wb_sm_35 (.D(n28767), .CK(clk), .Q(wb_sm)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(83[11] 90[18])
    defparam wb_sm_35.GSR = "ENABLED";
    LUT4 i13207_4_lut (.A(n29268), .B(wb_sm), .C(\address_7__N_549[1] ), 
         .D(spi_cmd_start), .Z(\address_7__N_565[1] )) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (B (C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(16[45:52])
    defparam i13207_4_lut.init = 16'he200;
    FD1P3AX wb_adr_i_i1 (.D(\address[1] ), .SP(wb_cyc_i_N_339), .CK(clk), 
            .Q(\wb_adr_i[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_adr_i_i1.GSR = "ENABLED";
    FD1P3AX wb_adr_i_i4 (.D(n29757), .SP(wb_cyc_i_N_339), .CK(clk), .Q(\wb_adr_i[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_adr_i_i4.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i1 (.D(wr_data[1]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i1.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i2 (.D(wr_data[2]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i2.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i3 (.D(wr_data[3]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i3.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i4 (.D(wr_data[4]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i4.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i5 (.D(wr_data[5]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i5.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i6 (.D(wr_data[6]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i6.GSR = "ENABLED";
    FD1P3AX wb_dat_i_i7 (.D(wr_data[7]), .SP(wb_we_i_N_344), .CK(clk), 
            .Q(wb_dat_i[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=15, LSE_LLINE=179, LSE_RLINE=196 */ ;   // c:/s_links/sources/wb_ctrl.v(101[11] 125[18])
    defparam wb_dat_i_i7.GSR = "ENABLED";
    LUT4 wr_en_I_0_1_lut (.A(wr_en), .Z(wr_en_N_355)) /* synthesis lut_function=(!(A)) */ ;   // c:/s_links/sources/wb_ctrl.v(129[44:50])
    defparam wr_en_I_0_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module spi_slave_efb
//

module spi_slave_efb (clk, n29239, wb_cyc_i, wb_we_i, GND_net, \wb_adr_i[4] , 
            \wb_adr_i[1] , \wb_adr_i[0] , wb_dat_i, spi_scsn_c, wb_dat_o, 
            \address_7__N_549[1] , spi_mosi_oe, spi_mosi_o, spi_miso_oe, 
            spi_miso_o, spi_clk_oe, spi_clk_o, spi_mosi_i, spi_miso_i, 
            spi_clk_i, VCC_net, n2720, mem_rdata_update_N_729, spi_addr_valid_N_732, 
            n29176, n2724, n29179, n7083, clk_enable_309, clk_enable_516, 
            wb_sm, clk_enable_95) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input clk;
    input n29239;
    input wb_cyc_i;
    input wb_we_i;
    input GND_net;
    input \wb_adr_i[4] ;
    input \wb_adr_i[1] ;
    input \wb_adr_i[0] ;
    input [7:0]wb_dat_i;
    input spi_scsn_c;
    output [7:0]wb_dat_o;
    output \address_7__N_549[1] ;
    output spi_mosi_oe;
    output spi_mosi_o;
    output spi_miso_oe;
    output spi_miso_o;
    output spi_clk_oe;
    output spi_clk_o;
    input spi_mosi_i;
    input spi_miso_i;
    input spi_clk_i;
    input VCC_net;
    input n2720;
    input mem_rdata_update_N_729;
    input spi_addr_valid_N_732;
    output n29176;
    input n2724;
    output n29179;
    input n7083;
    output clk_enable_309;
    output clk_enable_516;
    input wb_sm;
    output clk_enable_95;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire spi_clk_i /* synthesis is_clock=1 */ ;   // c:/s_links/sources/config_mcm/ip/spi_slave_efb.v(34[10:19])
    
    wire n29243;
    
    EFB EFBInst_0 (.WBCLKI(clk), .WBRSTI(n29239), .WBCYCI(wb_cyc_i), .WBSTBI(wb_cyc_i), 
        .WBWEI(wb_we_i), .WBADRI0(\wb_adr_i[0] ), .WBADRI1(\wb_adr_i[1] ), 
        .WBADRI2(GND_net), .WBADRI3(\wb_adr_i[4] ), .WBADRI4(\wb_adr_i[4] ), 
        .WBADRI5(GND_net), .WBADRI6(\wb_adr_i[4] ), .WBADRI7(GND_net), 
        .WBDATI0(wb_dat_i[0]), .WBDATI1(wb_dat_i[1]), .WBDATI2(wb_dat_i[2]), 
        .WBDATI3(wb_dat_i[3]), .WBDATI4(wb_dat_i[4]), .WBDATI5(wb_dat_i[5]), 
        .WBDATI6(wb_dat_i[6]), .WBDATI7(wb_dat_i[7]), .I2C1SCLI(GND_net), 
        .I2C1SDAI(GND_net), .I2C2SCLI(GND_net), .I2C2SDAI(GND_net), .SPISCKI(spi_clk_i), 
        .SPIMISOI(spi_miso_i), .SPIMOSII(spi_mosi_i), .SPISCSN(spi_scsn_c), 
        .TCCLKI(GND_net), .TCRSTN(GND_net), .TCIC(GND_net), .UFMSN(VCC_net), 
        .PLL0DATI0(GND_net), .PLL0DATI1(GND_net), .PLL0DATI2(GND_net), 
        .PLL0DATI3(GND_net), .PLL0DATI4(GND_net), .PLL0DATI5(GND_net), 
        .PLL0DATI6(GND_net), .PLL0DATI7(GND_net), .PLL0ACKI(GND_net), 
        .PLL1DATI0(GND_net), .PLL1DATI1(GND_net), .PLL1DATI2(GND_net), 
        .PLL1DATI3(GND_net), .PLL1DATI4(GND_net), .PLL1DATI5(GND_net), 
        .PLL1DATI6(GND_net), .PLL1DATI7(GND_net), .PLL1ACKI(GND_net), 
        .WBDATO0(wb_dat_o[0]), .WBDATO1(wb_dat_o[1]), .WBDATO2(wb_dat_o[2]), 
        .WBDATO3(wb_dat_o[3]), .WBDATO4(wb_dat_o[4]), .WBDATO5(wb_dat_o[5]), 
        .WBDATO6(wb_dat_o[6]), .WBDATO7(wb_dat_o[7]), .WBACKO(\address_7__N_549[1] ), 
        .SPISCKO(spi_clk_o), .SPISCKEN(spi_clk_oe), .SPIMISOO(spi_miso_o), 
        .SPIMISOEN(spi_miso_oe), .SPIMOSIO(spi_mosi_o), .SPIMOSIEN(spi_mosi_oe)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=6, LSE_LCOL=18, LSE_RCOL=15, LSE_LLINE=162, LSE_RLINE=176 */ ;   // c:/s_links/sources/spi_slave_top.v(162[18] 176[15])
    defparam EFBInst_0.EFB_I2C1 = "DISABLED";
    defparam EFBInst_0.EFB_I2C2 = "DISABLED";
    defparam EFBInst_0.EFB_SPI = "ENABLED";
    defparam EFBInst_0.EFB_TC = "DISABLED";
    defparam EFBInst_0.EFB_TC_PORTMODE = "WB";
    defparam EFBInst_0.EFB_UFM = "DISABLED";
    defparam EFBInst_0.EFB_WB_CLK_FREQ = "100.0";
    defparam EFBInst_0.DEV_DENSITY = "4000L";
    defparam EFBInst_0.UFM_INIT_PAGES = 0;
    defparam EFBInst_0.UFM_INIT_START_PAGE = 0;
    defparam EFBInst_0.UFM_INIT_ALL_ZEROS = "ENABLED";
    defparam EFBInst_0.UFM_INIT_FILE_NAME = "NONE";
    defparam EFBInst_0.UFM_INIT_FILE_FORMAT = "HEX";
    defparam EFBInst_0.I2C1_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C2_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C1_SLAVE_ADDR = "0b1000001";
    defparam EFBInst_0.I2C2_SLAVE_ADDR = "0b1000010";
    defparam EFBInst_0.I2C1_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C2_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C1_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C2_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C1_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C2_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C1_WAKEUP = "DISABLED";
    defparam EFBInst_0.I2C2_WAKEUP = "DISABLED";
    defparam EFBInst_0.SPI_MODE = "SLAVE";
    defparam EFBInst_0.SPI_CLK_DIVIDER = 2;
    defparam EFBInst_0.SPI_LSB_FIRST = "DISABLED";
    defparam EFBInst_0.SPI_CLK_INV = "DISABLED";
    defparam EFBInst_0.SPI_PHASE_ADJ = "DISABLED";
    defparam EFBInst_0.SPI_SLAVE_HANDSHAKE = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXOVR = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXOVR = "DISABLED";
    defparam EFBInst_0.SPI_WAKEUP = "DISABLED";
    defparam EFBInst_0.TC_MODE = "CTCM";
    defparam EFBInst_0.TC_SCLK_SEL = "PCLOCK";
    defparam EFBInst_0.TC_CCLK_SEL = 1;
    defparam EFBInst_0.GSR = "ENABLED";
    defparam EFBInst_0.TC_TOP_SET = 65535;
    defparam EFBInst_0.TC_OCR_SET = 32767;
    defparam EFBInst_0.TC_OC_MODE = "TOGGLE";
    defparam EFBInst_0.TC_RESETN = "ENABLED";
    defparam EFBInst_0.TC_TOP_SEL = "OFF";
    defparam EFBInst_0.TC_OV_INT = "OFF";
    defparam EFBInst_0.TC_OCR_INT = "OFF";
    defparam EFBInst_0.TC_ICR_INT = "OFF";
    defparam EFBInst_0.TC_OVERFLOW = "DISABLED";
    defparam EFBInst_0.TC_ICAPTURE = "DISABLED";
    LUT4 i72_2_lut_rep_515 (.A(n2720), .B(mem_rdata_update_N_729), .Z(n29243)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i72_2_lut_rep_515.init = 16'heeee;
    LUT4 i2_3_lut_rep_448_4_lut (.A(n2720), .B(mem_rdata_update_N_729), 
         .C(\address_7__N_549[1] ), .D(spi_addr_valid_N_732), .Z(n29176)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_3_lut_rep_448_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_451_3_lut (.A(n2720), .B(mem_rdata_update_N_729), 
         .C(n2724), .Z(n29179)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_rep_451_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n2720), .B(mem_rdata_update_N_729), .C(n7083), 
         .D(n2724), .Z(clk_enable_309)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i1_2_lut_4_lut (.A(spi_addr_valid_N_732), .B(n29243), .C(\address_7__N_549[1] ), 
         .D(n7083), .Z(clk_enable_516)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;   // c:/s_links/sources/spi_slave_top.v(162[18] 176[15])
    defparam i1_2_lut_4_lut.init = 16'hff20;
    LUT4 i22941_2_lut (.A(\address_7__N_549[1] ), .B(wb_sm), .Z(clk_enable_95)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/spi_slave_top.v(162[18] 176[15])
    defparam i22941_2_lut.init = 16'hbbbb;
    
endmodule
//
// Verilog Description of module spi_ctrl
//

module spi_ctrl (spi_addr_valid, clk, spi_addr_valid_N_732, clk_enable_516, 
            n29176, \address_7__N_549[1] , mem_rdata_update_N_729, resetn_c, 
            n29239, quad_set_complete, n29162, n29090, clk_enable_518, 
            spi_sdo_valid, clk_enable_523, n29127, n29211, n27225, 
            clk_enable_398, n29254, n29102, n29255, clk_enable_188, 
            n6, clk_enable_303, n32, \quad_homing[1] , n27657, n24, 
            n27201, n60, n29123, clk_enable_179, n29213, \spi_cmd_r[2] , 
            n29086, clk_enable_182, clear_intrpt, intrpt_out_N_2848, 
            n29100, clk_enable_185, wr_data, n29134, n27280, clk_enable_509, 
            reset_r_N_4813, EM_STOP, n29070, clk_enable_306, n29101, 
            \spi_addr_r[2] , clk_enable_186, quad_set_complete_adj_135, 
            n29120, clk_enable_505, \spi_addr_r[1] , n29111, clk_enable_76, 
            n29104, \spi_cmd_r[3] , clk_enable_436, n19233, clk_enable_184, 
            n29129, clk_enable_204, clear_intrpt_adj_136, intrpt_out_N_2635, 
            n29288, clk_enable_183, n29095, clk_enable_271, n29072, 
            n29083, clk_enable_521, quad_set_valid, n66, n21446, clk_1MHz_enable_171, 
            n29124, clk_enable_197, n26948, n13, n12714, n27301, 
            n29242, clk_enable_193, \spi_cmd_r[0] , n29074, clk_enable_200, 
            spi_sdo_valid_N_297, n10988, n29307, n27286, clk_enable_499, 
            n4, n27240, clk_enable_32, quad_set_complete_adj_137, n29092, 
            clk_enable_520, n29286, clk_enable_77, clear_intrpt_adj_138, 
            intrpt_out_N_2706, quad_set_valid_adj_139, n79, n20819, 
            clk_1MHz_enable_340, n27285, n29110, clk_enable_340, n31, 
            \quad_homing[1]_adj_140 , n5, n26, n27234, clk_enable_174, 
            n27243, clk_enable_171, clk_enable_172, n29119, n29174, 
            clk_enable_435, n29082, n29106, clk_enable_506, \spi_data[0] , 
            wb_dat_o, n29144, clk_enable_269, n13074, clk_enable_167, 
            n29175, clk_enable_28, clk_enable_309, n29179, n27259, 
            n29107, clk_enable_131, clear_intrpt_adj_141, intrpt_out_N_2919, 
            n65, clk_enable_194, n65_adj_142, clk_enable_177, spi_sdo_valid_N_296, 
            clk_enable_305, clk_enable_189, \address[0] , clk_enable_180, 
            wr_en, spi_scsn_c, clk_enable_162, clk_enable_166, n29256, 
            clk_enable_175, clk_enable_176, quad_set_complete_adj_143, 
            n29105, clk_enable_502, n29071, n29077, clk_enable_526, 
            n29069, n29075, clk_enable_342, clk_enable_202, clear_intrpt_adj_144, 
            intrpt_out_N_2990, clk_enable_201, clk_enable_467, clk_enable_191, 
            clk_enable_187, clk_enable_192, quad_set_complete_adj_145, 
            clk_enable_519, clk_enable_170, n29118, n29214, clk_enable_286, 
            n29182, clk_enable_359, reset_r_N_4474, n29097, clk_enable_307, 
            clear_intrpt_adj_146, intrpt_out_N_3061, clk_enable_86, clk_enable_181, 
            clk_enable_288, clk_enable_433, clk_enable_434, quad_set_complete_adj_147, 
            clk_enable_501, n29205, clk_enable_169, clear_intrpt_adj_148, 
            intrpt_out_N_2777, n27058, clk_enable_400, clk_enable_402, 
            quad_set_complete_adj_149, clk_enable_503, clk_enable_30, 
            n2724, n2720, spi_cmd, wr_en_N_355, n9633, spi_addr, 
            n27465, n26928, n29141, n29126, n27618, spi_cmd_start, 
            n29268, wb_sm, n28767, wb_cyc_i_N_339, \address_7__N_565[1] , 
            n7083, mem_rdata, GND_net, n29114, clk_enable_20, \spi_data[1] , 
            \spi_data[2] , \spi_data[3] , \spi_data[4] , \spi_data[5] , 
            \spi_data[6] , \spi_data[7] , \spi_data[8] , \spi_data[9] , 
            \spi_data[10] , \spi_data[11] , \spi_data[12] , \spi_data[13] , 
            \spi_data[14] , \spi_data[15] , \spi_data[16] , \spi_data[17] , 
            \spi_data[18] , \spi_data[19] , \spi_data[20] , \spi_data[21] , 
            \spi_data[22] , \spi_data[23] , \spi_data[24] , \spi_data[25] , 
            \spi_data[26] , \spi_data[27] , \spi_data[28] , \spi_data[29] , 
            \spi_data[30] , \spi_data[31] , \address[1] , spi_data_valid, 
            spi_cmd_valid, n31_adj_150, wb_we_i_N_344, n29761) /* synthesis syn_module_defined=1 */ ;
    output spi_addr_valid;
    input clk;
    output spi_addr_valid_N_732;
    input clk_enable_516;
    input n29176;
    input \address_7__N_549[1] ;
    output mem_rdata_update_N_729;
    input resetn_c;
    output n29239;
    input quad_set_complete;
    input n29162;
    input n29090;
    output clk_enable_518;
    input spi_sdo_valid;
    output clk_enable_523;
    input n29127;
    input n29211;
    input n27225;
    output clk_enable_398;
    input n29254;
    input n29102;
    input n29255;
    output clk_enable_188;
    input n6;
    output clk_enable_303;
    input n32;
    input \quad_homing[1] ;
    input n27657;
    output n24;
    input n27201;
    input n60;
    input n29123;
    output clk_enable_179;
    input n29213;
    input \spi_cmd_r[2] ;
    input n29086;
    output clk_enable_182;
    input clear_intrpt;
    output intrpt_out_N_2848;
    input n29100;
    output clk_enable_185;
    output [7:0]wr_data;
    input n29134;
    input n27280;
    output clk_enable_509;
    input reset_r_N_4813;
    input EM_STOP;
    input n29070;
    output clk_enable_306;
    input n29101;
    input \spi_addr_r[2] ;
    output clk_enable_186;
    input quad_set_complete_adj_135;
    input n29120;
    output clk_enable_505;
    input \spi_addr_r[1] ;
    input n29111;
    output clk_enable_76;
    input n29104;
    input \spi_cmd_r[3] ;
    output clk_enable_436;
    input n19233;
    output clk_enable_184;
    input n29129;
    output clk_enable_204;
    input clear_intrpt_adj_136;
    output intrpt_out_N_2635;
    input n29288;
    output clk_enable_183;
    input n29095;
    output clk_enable_271;
    input n29072;
    input n29083;
    output clk_enable_521;
    input quad_set_valid;
    input n66;
    input n21446;
    output clk_1MHz_enable_171;
    input n29124;
    output clk_enable_197;
    input n26948;
    input n13;
    input n12714;
    output n27301;
    input n29242;
    output clk_enable_193;
    input \spi_cmd_r[0] ;
    input n29074;
    output clk_enable_200;
    input spi_sdo_valid_N_297;
    output n10988;
    input n29307;
    input n27286;
    output clk_enable_499;
    input n4;
    input n27240;
    output clk_enable_32;
    input quad_set_complete_adj_137;
    input n29092;
    output clk_enable_520;
    input n29286;
    output clk_enable_77;
    input clear_intrpt_adj_138;
    output intrpt_out_N_2706;
    input quad_set_valid_adj_139;
    input n79;
    input n20819;
    output clk_1MHz_enable_340;
    input n27285;
    input n29110;
    output clk_enable_340;
    input n31;
    input \quad_homing[1]_adj_140 ;
    input n5;
    output n26;
    input n27234;
    output clk_enable_174;
    input n27243;
    output clk_enable_171;
    output clk_enable_172;
    input n29119;
    input n29174;
    output clk_enable_435;
    input n29082;
    input n29106;
    output clk_enable_506;
    output \spi_data[0] ;
    input [7:0]wb_dat_o;
    input n29144;
    output clk_enable_269;
    input n13074;
    output clk_enable_167;
    input n29175;
    output clk_enable_28;
    input clk_enable_309;
    input n29179;
    input n27259;
    input n29107;
    output clk_enable_131;
    input clear_intrpt_adj_141;
    output intrpt_out_N_2919;
    input n65;
    output clk_enable_194;
    input n65_adj_142;
    output clk_enable_177;
    input spi_sdo_valid_N_296;
    output clk_enable_305;
    output clk_enable_189;
    output \address[0] ;
    output clk_enable_180;
    output wr_en;
    input spi_scsn_c;
    output clk_enable_162;
    output clk_enable_166;
    input n29256;
    output clk_enable_175;
    output clk_enable_176;
    input quad_set_complete_adj_143;
    input n29105;
    output clk_enable_502;
    input n29071;
    input n29077;
    output clk_enable_526;
    input n29069;
    input n29075;
    output clk_enable_342;
    output clk_enable_202;
    input clear_intrpt_adj_144;
    output intrpt_out_N_2990;
    output clk_enable_201;
    output clk_enable_467;
    output clk_enable_191;
    output clk_enable_187;
    output clk_enable_192;
    input quad_set_complete_adj_145;
    output clk_enable_519;
    output clk_enable_170;
    input n29118;
    input n29214;
    output clk_enable_286;
    input n29182;
    output clk_enable_359;
    input reset_r_N_4474;
    input n29097;
    output clk_enable_307;
    input clear_intrpt_adj_146;
    output intrpt_out_N_3061;
    output clk_enable_86;
    output clk_enable_181;
    output clk_enable_288;
    output clk_enable_433;
    output clk_enable_434;
    input quad_set_complete_adj_147;
    output clk_enable_501;
    input n29205;
    output clk_enable_169;
    input clear_intrpt_adj_148;
    output intrpt_out_N_2777;
    input n27058;
    output clk_enable_400;
    output clk_enable_402;
    input quad_set_complete_adj_149;
    output clk_enable_503;
    output clk_enable_30;
    output n2724;
    output n2720;
    output [15:0]spi_cmd;
    input wr_en_N_355;
    input n9633;
    output [7:0]spi_addr;
    output n27465;
    output n26928;
    output n29141;
    output n29126;
    output n27618;
    output spi_cmd_start;
    output n29268;
    input wb_sm;
    output n28767;
    output wb_cyc_i_N_339;
    input \address_7__N_565[1] ;
    output n7083;
    input [7:0]mem_rdata;
    input GND_net;
    input n29114;
    output clk_enable_20;
    output \spi_data[1] ;
    output \spi_data[2] ;
    output \spi_data[3] ;
    output \spi_data[4] ;
    output \spi_data[5] ;
    output \spi_data[6] ;
    output \spi_data[7] ;
    output \spi_data[8] ;
    output \spi_data[9] ;
    output \spi_data[10] ;
    output \spi_data[11] ;
    output \spi_data[12] ;
    output \spi_data[13] ;
    output \spi_data[14] ;
    output \spi_data[15] ;
    output \spi_data[16] ;
    output \spi_data[17] ;
    output \spi_data[18] ;
    output \spi_data[19] ;
    output \spi_data[20] ;
    output \spi_data[21] ;
    output \spi_data[22] ;
    output \spi_data[23] ;
    output \spi_data[24] ;
    output \spi_data[25] ;
    output \spi_data[26] ;
    output \spi_data[27] ;
    output \spi_data[28] ;
    output \spi_data[29] ;
    output \spi_data[30] ;
    output \spi_data[31] ;
    output \address[1] ;
    output spi_data_valid;
    output spi_cmd_valid;
    output n31_adj_150;
    output wb_we_i_N_344;
    output n29761;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    wire clk_enable_3;
    wire [3:0]spi_byte_cnt;   // c:/s_links/sources/spi_ctrl.v(74[13:25])
    wire [3:0]n21;
    
    wire n29308;
    wire [15:0]n2713;
    
    wire n29238, n29173, mem_rdata_update, clk_enable_366;
    wire [7:0]n672;
    
    wire spi_cmd_start_reg_N_745, n26429, n28855, n28854, n29186, 
        n28856, clk_enable_474, n7710;
    wire [7:0]mem_burst_cnt;   // c:/s_links/sources/spi_ctrl.v(71[16:29])
    wire [7:0]n37;
    
    wire spi_idle_N_747, spi_csn_buf0_p, spi_csn_buf2_p, spi_cmd_start_reg, 
        n28766, spi_idle, n14197;
    wire [7:0]address_7__N_359;
    
    wire rd_en, rd_en_N_710, wr_en_N_697, spi_cmd_cnt, spi_cmd_cnt_N_749, 
        spi_cmd_start_reg_N_746, n29240, n4606, n29241, n29318, n5876, 
        n29248, n10729, n29073, n29252, n29180, n29269, n26_adj_6703, 
        n38_adj_6704, n9972, n19324, n27601, n28765, n28764;
    wire [7:0]n47;
    
    wire n29262, n22_adj_6705, n8, n5874, n5880;
    wire [1:0]n6901;
    
    wire n27679, n29266, n29136, n4_adj_6706, wr_en_N_703, n29143, 
        n29142, n27180, n29319, n27578, n29187, clk_enable_504, 
        n27630, spi_data_valid_N_737, n26945, clk_enable_482, n10, 
        clk_enable_490, clk_enable_498, n28722, n29128, n29125, rd_en_N_717, 
        n4_adj_6707, n25453, n32_adj_6708, n27675, n29279, clk_enable_525, 
        clk_enable_279;
    wire [7:0]n37_adj_6725;
    
    wire n8_adj_6709, mem_wr_N_726, n19198, n26923, n25199, n25198, 
        n25197, n25196, n25195, n25194, n25193, n25192, n18948, 
        clk_enable_507, n36, n28723, n18, n15, n13622, n30, n9429, 
        n26319, n9988, n9986, n25364, n9982, n9980, n9976, n13_adj_6718, 
        n18908, mem_wr, n2775, n6_adj_6720, n29116, n4_adj_6721, 
        n4_adj_6722, n10_adj_6723, n12, n4_adj_6724, n13568, n27596, 
        n13657, n7;
    
    FD1P3AX spi_addr_valid_224 (.D(spi_addr_valid_N_732), .SP(clk_enable_3), 
            .CK(clk), .Q(spi_addr_valid)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_addr_valid_224.GSR = "ENABLED";
    FD1P3IX spi_byte_cnt_2505__i3 (.D(n21[3]), .SP(clk_enable_516), .CD(n29176), 
            .CK(clk), .Q(spi_byte_cnt[3]));   // c:/s_links/sources/spi_ctrl.v(383[46:62])
    defparam spi_byte_cnt_2505__i3.GSR = "ENABLED";
    FD1P3IX spi_byte_cnt_2505__i2 (.D(n21[2]), .SP(clk_enable_516), .CD(n29176), 
            .CK(clk), .Q(spi_byte_cnt[2]));   // c:/s_links/sources/spi_ctrl.v(383[46:62])
    defparam spi_byte_cnt_2505__i2.GSR = "ENABLED";
    LUT4 i15_4_lut (.A(n29308), .B(\address_7__N_549[1] ), .C(spi_addr_valid_N_732), 
         .D(n2713[11]), .Z(clk_enable_3)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(16[45:52])
    defparam i15_4_lut.init = 16'hcfca;
    LUT4 i2_3_lut_rep_510 (.A(n2713[6]), .B(n2713[2]), .C(mem_rdata_update_N_729), 
         .Z(n29238)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i2_3_lut_rep_510.init = 16'hfefe;
    LUT4 i1_2_lut_rep_445_4_lut (.A(n2713[6]), .B(n2713[2]), .C(mem_rdata_update_N_729), 
         .D(spi_addr_valid_N_732), .Z(n29173)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_2_lut_rep_445_4_lut.init = 16'hfffe;
    LUT4 resetn_I_0_1_lut_rep_511 (.A(resetn_c), .Z(n29239)) /* synthesis lut_function=(!(A)) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_I_0_1_lut_rep_511.init = 16'h5555;
    LUT4 i2_3_lut_4_lut_4_lut (.A(resetn_c), .B(quad_set_complete), .C(n29162), 
         .D(n29090), .Z(clk_enable_518)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_3_lut_4_lut_4_lut.init = 16'hfddd;
    LUT4 i2_3_lut_3_lut (.A(resetn_c), .B(mem_rdata_update), .C(spi_sdo_valid), 
         .Z(clk_enable_523)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_3_lut_3_lut.init = 16'hfdfd;
    LUT4 i2745_2_lut_4_lut_4_lut (.A(resetn_c), .B(n29127), .C(n29211), 
         .D(n27225), .Z(clk_enable_398)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2745_2_lut_4_lut_4_lut.init = 16'hd555;
    LUT4 i1_3_lut_4_lut_4_lut (.A(resetn_c), .B(n29254), .C(n29102), .D(n29255), 
         .Z(clk_enable_188)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 i2735_2_lut_2_lut (.A(resetn_c), .B(n6), .Z(clk_enable_303)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2735_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_4_lut_4_lut (.A(resetn_c), .B(n32), .C(\quad_homing[1] ), 
         .D(n27657), .Z(n24)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_4_lut.init = 16'h5d55;
    LUT4 i2919_3_lut_4_lut_4_lut (.A(resetn_c), .B(n27201), .C(n60), .D(n29123), 
         .Z(clk_enable_179)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2919_3_lut_4_lut_4_lut.init = 16'hd555;
    LUT4 i1_4_lut_4_lut_adj_483 (.A(resetn_c), .B(n29213), .C(\spi_cmd_r[2] ), 
         .D(n29086), .Z(clk_enable_182)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_4_lut_adj_483.init = 16'hd555;
    LUT4 resetn_N_2845_I_0_2_lut_2_lut (.A(resetn_c), .B(clear_intrpt), 
         .Z(intrpt_out_N_2848)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_N_2845_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i2967_3_lut_4_lut_4_lut (.A(resetn_c), .B(n29254), .C(n29100), 
         .D(n29255), .Z(clk_enable_185)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2967_3_lut_4_lut_4_lut.init = 16'h55d5;
    FD1P3AX wr_data_i0_i0 (.D(n672[0]), .SP(clk_enable_366), .CK(clk), 
            .Q(wr_data[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i0.GSR = "ENABLED";
    LUT4 i2737_4_lut_4_lut (.A(resetn_c), .B(n29134), .C(\spi_cmd_r[2] ), 
         .D(n27280), .Z(clk_enable_509)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2737_4_lut_4_lut.init = 16'hd555;
    LUT4 i2_4_lut_4_lut (.A(resetn_c), .B(reset_r_N_4813), .C(EM_STOP), 
         .D(n29070), .Z(clk_enable_306)) /* synthesis lut_function=((B (D)+!B (C+(D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_4_lut_4_lut.init = 16'hff75;
    LUT4 i1_3_lut_4_lut_4_lut_adj_484 (.A(resetn_c), .B(\spi_cmd_r[2] ), 
         .C(n29101), .D(\spi_addr_r[2] ), .Z(clk_enable_186)) /* synthesis lut_function=(!(A (B+((D)+!C)))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_484.init = 16'h5575;
    LUT4 i2_3_lut_3_lut_adj_485 (.A(resetn_c), .B(quad_set_complete_adj_135), 
         .C(n29120), .Z(clk_enable_505)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_3_lut_3_lut_adj_485.init = 16'hfdfd;
    LUT4 i1_2_lut_4_lut_4_lut (.A(resetn_c), .B(n29162), .C(\spi_addr_r[1] ), 
         .D(n29111), .Z(clk_enable_76)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_4_lut_4_lut.init = 16'hd555;
    LUT4 i2738_3_lut_3_lut (.A(resetn_c), .B(n29104), .C(\spi_cmd_r[3] ), 
         .Z(clk_enable_436)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2738_3_lut_3_lut.init = 16'h5d5d;
    LUT4 i2861_3_lut_4_lut_4_lut (.A(resetn_c), .B(n27201), .C(n29123), 
         .D(n19233), .Z(clk_enable_184)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2861_3_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 i2947_4_lut_4_lut (.A(resetn_c), .B(n29213), .C(n29129), .D(n27225), 
         .Z(clk_enable_204)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2947_4_lut_4_lut.init = 16'hd555;
    FD1P3IX spi_byte_cnt_2505__i1 (.D(n21[1]), .SP(clk_enable_516), .CD(n29176), 
            .CK(clk), .Q(spi_byte_cnt[1]));   // c:/s_links/sources/spi_ctrl.v(383[46:62])
    defparam spi_byte_cnt_2505__i1.GSR = "ENABLED";
    LUT4 resetn_N_2632_I_0_2_lut_2_lut (.A(resetn_c), .B(clear_intrpt_adj_136), 
         .Z(intrpt_out_N_2635)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_N_2632_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_4_lut_4_lut_adj_486 (.A(resetn_c), .B(n29288), .C(n29254), 
         .D(n29100), .Z(clk_enable_183)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_4_lut_adj_486.init = 16'hd555;
    LUT4 i2789_2_lut_3_lut_4_lut_4_lut (.A(resetn_c), .B(n29255), .C(n29095), 
         .D(\spi_cmd_r[2] ), .Z(clk_enable_271)) /* synthesis lut_function=(!(A (B+((D)+!C)))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2789_2_lut_3_lut_4_lut_4_lut.init = 16'h5575;
    FD1S3AY main_sm_FSM_i1 (.D(n26429), .CK(clk), .Q(spi_cmd_start_reg_N_745));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i1.GSR = "ENABLED";
    LUT4 i2_4_lut_4_lut_adj_487 (.A(resetn_c), .B(EM_STOP), .C(n29072), 
         .D(n29083), .Z(clk_enable_521)) /* synthesis lut_function=((B ((D)+!C)+!B (D))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_4_lut_4_lut_adj_487.init = 16'hff5d;
    LUT4 i2_4_lut_4_lut_adj_488 (.A(resetn_c), .B(quad_set_valid), .C(n66), 
         .D(n21446), .Z(clk_1MHz_enable_171)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_4_lut_4_lut_adj_488.init = 16'hfffd;
    LUT4 i1_3_lut_4_lut_4_lut_adj_489 (.A(resetn_c), .B(n29213), .C(n29124), 
         .D(n29129), .Z(clk_enable_197)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_489.init = 16'h5d55;
    LUT4 i1_4_lut_4_lut_adj_490 (.A(resetn_c), .B(n26948), .C(n13), .D(n12714), 
         .Z(n27301)) /* synthesis lut_function=((B (D)+!B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_4_lut_adj_490.init = 16'hfd55;
    LUT4 i2951_3_lut_4_lut_4_lut (.A(resetn_c), .B(n29242), .C(n29095), 
         .D(\spi_cmd_r[2] ), .Z(clk_enable_193)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2951_3_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 i2943_4_lut_4_lut (.A(resetn_c), .B(\spi_cmd_r[0] ), .C(n29255), 
         .D(n29074), .Z(clk_enable_200)) /* synthesis lut_function=(!(A (B+(C+!(D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2943_4_lut_4_lut.init = 16'h5755;
    LUT4 i6188_2_lut_2_lut (.A(resetn_c), .B(spi_sdo_valid_N_297), .Z(n10988)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i6188_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_3_lut_4_lut_4_lut_adj_491 (.A(resetn_c), .B(n29307), .C(n27286), 
         .D(n29111), .Z(clk_enable_499)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_491.init = 16'hd555;
    LUT4 i1_3_lut_4_lut_4_lut_adj_492 (.A(resetn_c), .B(n4), .C(n27240), 
         .D(n29123), .Z(clk_enable_32)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_492.init = 16'hd555;
    LUT4 i2_3_lut_3_lut_adj_493 (.A(resetn_c), .B(quad_set_complete_adj_137), 
         .C(n29092), .Z(clk_enable_520)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_3_lut_3_lut_adj_493.init = 16'hfdfd;
    PFUMX i23093 (.BLUT(n28855), .ALUT(n28854), .C0(n29186), .Z(n28856));
    LUT4 i1_3_lut_4_lut_4_lut_adj_494 (.A(resetn_c), .B(n29286), .C(n27286), 
         .D(n29111), .Z(clk_enable_77)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_494.init = 16'h7555;
    LUT4 resetn_N_2703_I_0_2_lut_2_lut (.A(resetn_c), .B(clear_intrpt_adj_138), 
         .Z(intrpt_out_N_2706)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_N_2703_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i2_4_lut_4_lut_adj_495 (.A(resetn_c), .B(quad_set_valid_adj_139), 
         .C(n79), .D(n20819), .Z(clk_1MHz_enable_340)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_4_lut_4_lut_adj_495.init = 16'hfffd;
    LUT4 i2_4_lut_4_lut_adj_496 (.A(resetn_c), .B(EM_STOP), .C(n27285), 
         .D(n29110), .Z(clk_enable_340)) /* synthesis lut_function=((B ((D)+!C)+!B (D))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_4_lut_4_lut_adj_496.init = 16'hff5d;
    LUT4 i1_4_lut_4_lut_adj_497 (.A(resetn_c), .B(n31), .C(\quad_homing[1]_adj_140 ), 
         .D(n5), .Z(n26)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_4_lut_4_lut_adj_497.init = 16'h5d55;
    LUT4 i2979_3_lut_3_lut (.A(resetn_c), .B(n27234), .C(\spi_addr_r[2] ), 
         .Z(clk_enable_174)) /* synthesis lut_function=((B (C))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2979_3_lut_3_lut.init = 16'hd5d5;
    LUT4 i2927_3_lut_4_lut_4_lut (.A(resetn_c), .B(n27243), .C(n60), .D(n29123), 
         .Z(clk_enable_171)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2927_3_lut_4_lut_4_lut.init = 16'hd555;
    LUT4 i2935_3_lut_4_lut_4_lut (.A(resetn_c), .B(n29211), .C(n29086), 
         .D(\spi_cmd_r[2] ), .Z(clk_enable_172)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2935_3_lut_4_lut_4_lut.init = 16'hd555;
    LUT4 i2742_4_lut_4_lut (.A(resetn_c), .B(n29119), .C(n29174), .D(n27240), 
         .Z(clk_enable_435)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2742_4_lut_4_lut.init = 16'hd555;
    LUT4 i2_4_lut_4_lut_adj_498 (.A(resetn_c), .B(n29082), .C(EM_STOP), 
         .D(n29106), .Z(clk_enable_506)) /* synthesis lut_function=((B (D)+!B (C+(D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_4_lut_4_lut_adj_498.init = 16'hff75;
    FD1P3IX spi_data__i0 (.D(wb_dat_o[0]), .SP(clk_enable_474), .CD(n7710), 
            .CK(clk), .Q(\spi_data[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i0.GSR = "ENABLED";
    LUT4 i2743_2_lut_3_lut_4_lut_4_lut (.A(resetn_c), .B(n29134), .C(n29144), 
         .D(\spi_cmd_r[2] ), .Z(clk_enable_269)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2743_2_lut_3_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 i1_3_lut_4_lut_4_lut_adj_499 (.A(resetn_c), .B(n13074), .C(n29124), 
         .D(n29129), .Z(clk_enable_167)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_499.init = 16'h5d55;
    LUT4 i2748_3_lut_4_lut_4_lut (.A(resetn_c), .B(n29175), .C(n29090), 
         .D(n29174), .Z(clk_enable_28)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2748_3_lut_4_lut_4_lut.init = 16'hd555;
    FD1P3IX mem_burst_cnt_2507__i7 (.D(n37[7]), .SP(clk_enable_309), .CD(n29179), 
            .CK(clk), .Q(mem_burst_cnt[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_2507__i7.GSR = "ENABLED";
    FD1P3IX mem_burst_cnt_2507__i6 (.D(n37[6]), .SP(clk_enable_309), .CD(n29179), 
            .CK(clk), .Q(mem_burst_cnt[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_2507__i6.GSR = "ENABLED";
    FD1S3AY spi_csn_buf1_p_209 (.D(spi_csn_buf0_p), .CK(clk), .Q(spi_idle_N_747)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(103[11:44])
    defparam spi_csn_buf1_p_209.GSR = "ENABLED";
    FD1S3AY spi_csn_buf2_p_210 (.D(spi_idle_N_747), .CK(clk), .Q(spi_csn_buf2_p)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(110[11:44])
    defparam spi_csn_buf2_p_210.GSR = "ENABLED";
    FD1S3AX spi_cmd_start_reg_211 (.D(n28766), .CK(clk), .Q(spi_cmd_start_reg)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(117[11] 120[40])
    defparam spi_cmd_start_reg_211.GSR = "ENABLED";
    FD1S3AX spi_idle_212 (.D(n14197), .CK(clk), .Q(spi_idle)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(130[11] 133[31])
    defparam spi_idle_212.GSR = "ENABLED";
    FD1P3IX mem_burst_cnt_2507__i5 (.D(n37[5]), .SP(clk_enable_309), .CD(n29179), 
            .CK(clk), .Q(mem_burst_cnt[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_2507__i5.GSR = "ENABLED";
    FD1P3IX mem_burst_cnt_2507__i4 (.D(n37[4]), .SP(clk_enable_309), .CD(n29179), 
            .CK(clk), .Q(mem_burst_cnt[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_2507__i4.GSR = "ENABLED";
    FD1P3IX mem_burst_cnt_2507__i3 (.D(n37[3]), .SP(clk_enable_309), .CD(n29179), 
            .CK(clk), .Q(mem_burst_cnt[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_2507__i3.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(resetn_c), .B(n27259), .C(n29107), 
         .D(\spi_cmd_r[2] ), .Z(clk_enable_131)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 resetn_N_2916_I_0_2_lut_2_lut (.A(resetn_c), .B(clear_intrpt_adj_141), 
         .Z(intrpt_out_N_2919)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_N_2916_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i2955_4_lut_4_lut (.A(resetn_c), .B(n4), .C(n29242), .D(n65), 
         .Z(clk_enable_194)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2955_4_lut_4_lut.init = 16'hd555;
    LUT4 i2975_3_lut_4_lut_4_lut (.A(resetn_c), .B(n65_adj_142), .C(n29102), 
         .D(n29255), .Z(clk_enable_177)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2975_3_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 i1_2_lut_2_lut (.A(resetn_c), .B(spi_sdo_valid_N_296), .Z(clk_enable_305)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_2_lut.init = 16'hdddd;
    LUT4 i2915_3_lut_4_lut_4_lut (.A(resetn_c), .B(\spi_cmd_r[2] ), .C(n29101), 
         .D(\spi_addr_r[2] ), .Z(clk_enable_189)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2915_3_lut_4_lut_4_lut.init = 16'h55d5;
    FD1S3AY address_i1 (.D(address_7__N_359[0]), .CK(clk), .Q(\address[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam address_i1.GSR = "ENABLED";
    LUT4 i2869_3_lut_4_lut_4_lut (.A(resetn_c), .B(n27243), .C(n29123), 
         .D(n19233), .Z(clk_enable_180)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2869_3_lut_4_lut_4_lut.init = 16'h55d5;
    FD1S3AX rd_en_215 (.D(rd_en_N_710), .CK(clk), .Q(rd_en)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam rd_en_215.GSR = "ENABLED";
    FD1S3AX wr_en_216 (.D(wr_en_N_697), .CK(clk), .Q(wr_en)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_en_216.GSR = "ENABLED";
    FD1S3AX spi_cmd_cnt_228 (.D(spi_cmd_cnt_N_749), .CK(clk), .Q(spi_cmd_cnt)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_cnt_228.GSR = "ENABLED";
    FD1S3AY spi_csn_buf0_p_208 (.D(spi_scsn_c), .CK(clk), .Q(spi_csn_buf0_p)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(96[11:37])
    defparam spi_csn_buf0_p_208.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_500 (.A(resetn_c), .B(n29162), .C(n29107), 
         .D(\spi_cmd_r[2] ), .Z(clk_enable_162)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_500.init = 16'h55d5;
    LUT4 i1_3_lut_4_lut_4_lut_adj_501 (.A(resetn_c), .B(n13074), .C(n29086), 
         .D(\spi_cmd_r[2] ), .Z(clk_enable_166)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_501.init = 16'hd555;
    LUT4 i2879_3_lut_4_lut_4_lut (.A(resetn_c), .B(n27201), .C(n29256), 
         .D(n29123), .Z(clk_enable_175)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2879_3_lut_4_lut_4_lut.init = 16'hd555;
    LUT4 i1_3_lut_4_lut_4_lut_adj_502 (.A(resetn_c), .B(n60), .C(n27240), 
         .D(n29123), .Z(clk_enable_176)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_502.init = 16'hd555;
    LUT4 i2_3_lut_4_lut_4_lut_adj_503 (.A(resetn_c), .B(quad_set_complete_adj_143), 
         .C(n27259), .D(n29105), .Z(clk_enable_502)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_3_lut_4_lut_4_lut_adj_503.init = 16'hfddd;
    LUT4 i2_4_lut_4_lut_adj_504 (.A(resetn_c), .B(n29071), .C(EM_STOP), 
         .D(n29077), .Z(clk_enable_526)) /* synthesis lut_function=((B (D)+!B (C+(D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_4_lut_4_lut_adj_504.init = 16'hff75;
    LUT4 i2_4_lut_4_lut_adj_505 (.A(resetn_c), .B(n29069), .C(EM_STOP), 
         .D(n29075), .Z(clk_enable_342)) /* synthesis lut_function=((B (D)+!B (C+(D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_4_lut_4_lut_adj_505.init = 16'hff75;
    LUT4 i1_3_lut_4_lut_4_lut_adj_506 (.A(resetn_c), .B(n29255), .C(n29095), 
         .D(\spi_cmd_r[2] ), .Z(clk_enable_202)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_506.init = 16'h7555;
    LUT4 resetn_N_2987_I_0_2_lut_2_lut (.A(resetn_c), .B(clear_intrpt_adj_144), 
         .Z(intrpt_out_N_2990)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_N_2987_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_3_lut_4_lut_4_lut_adj_507 (.A(resetn_c), .B(n29288), .C(n29095), 
         .D(\spi_cmd_r[2] ), .Z(clk_enable_201)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_507.init = 16'hd555;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_508 (.A(resetn_c), .B(n27259), .C(n29119), 
         .D(\spi_addr_r[1] ), .Z(clk_enable_467)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_508.init = 16'h55d5;
    LUT4 i2911_3_lut_4_lut_4_lut (.A(resetn_c), .B(n4), .C(n65), .D(n29255), 
         .Z(clk_enable_191)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2911_3_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 i2963_3_lut_3_lut (.A(resetn_c), .B(n27234), .C(\spi_addr_r[2] ), 
         .Z(clk_enable_187)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2963_3_lut_3_lut.init = 16'h5d5d;
    LUT4 i2959_3_lut_4_lut_4_lut (.A(resetn_c), .B(n65_adj_142), .C(n29100), 
         .D(n29255), .Z(clk_enable_192)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2959_3_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 i2_3_lut_4_lut_4_lut_adj_509 (.A(resetn_c), .B(quad_set_complete_adj_145), 
         .C(n27259), .D(n29090), .Z(clk_enable_519)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_3_lut_4_lut_4_lut_adj_509.init = 16'hfddd;
    LUT4 i1_3_lut_4_lut_4_lut_adj_510 (.A(resetn_c), .B(n29256), .C(n27240), 
         .D(n29123), .Z(clk_enable_170)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_510.init = 16'hd555;
    LUT4 i1_3_lut_4_lut_4_lut_adj_511 (.A(resetn_c), .B(n27201), .C(n29118), 
         .D(n29214), .Z(clk_enable_286)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_511.init = 16'h55d5;
    LUT4 i1_2_lut_4_lut_4_lut_adj_512 (.A(resetn_c), .B(n29182), .C(n29090), 
         .D(n13074), .Z(clk_enable_359)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_4_lut_4_lut_adj_512.init = 16'h7555;
    LUT4 i2_4_lut_4_lut_adj_513 (.A(resetn_c), .B(reset_r_N_4474), .C(EM_STOP), 
         .D(n29097), .Z(clk_enable_307)) /* synthesis lut_function=((B (D)+!B (C+(D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_4_lut_4_lut_adj_513.init = 16'hff75;
    LUT4 resetn_N_3058_I_0_2_lut_2_lut (.A(resetn_c), .B(clear_intrpt_adj_146), 
         .Z(intrpt_out_N_3061)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_N_3058_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_4_lut_4_lut_adj_514 (.A(resetn_c), .B(n65), .C(n29288), 
         .D(n19233), .Z(clk_enable_86)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_4_lut_4_lut_adj_514.init = 16'h55d5;
    LUT4 i1_3_lut_4_lut_4_lut_adj_515 (.A(resetn_c), .B(n19233), .C(n27240), 
         .D(n29123), .Z(clk_enable_181)) /* synthesis lut_function=(!(A (B+!(C (D))))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_515.init = 16'h7555;
    LUT4 i2849_2_lut_3_lut_4_lut_4_lut (.A(resetn_c), .B(n29256), .C(n65), 
         .D(n29255), .Z(clk_enable_288)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2849_2_lut_3_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_516 (.A(resetn_c), .B(n29162), .C(n29119), 
         .D(\spi_addr_r[1] ), .Z(clk_enable_433)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_516.init = 16'h55d5;
    LUT4 i1_3_lut_4_lut_4_lut_adj_517 (.A(resetn_c), .B(n27243), .C(n29118), 
         .D(n29214), .Z(clk_enable_434)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_517.init = 16'h55d5;
    LUT4 i2_3_lut_4_lut_4_lut_adj_518 (.A(resetn_c), .B(quad_set_complete_adj_147), 
         .C(n29105), .D(n29162), .Z(clk_enable_501)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_3_lut_4_lut_4_lut_adj_518.init = 16'hfddd;
    LUT4 i1_3_lut_4_lut_4_lut_adj_519 (.A(resetn_c), .B(n29205), .C(n29086), 
         .D(\spi_cmd_r[2] ), .Z(clk_enable_169)) /* synthesis lut_function=((B (C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_3_lut_4_lut_4_lut_adj_519.init = 16'hd555;
    LUT4 resetn_N_2774_I_0_2_lut_2_lut (.A(resetn_c), .B(clear_intrpt_adj_148), 
         .Z(intrpt_out_N_2777)) /* synthesis lut_function=((B)+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam resetn_N_2774_I_0_2_lut_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_520 (.A(resetn_c), .B(n27058), .C(n29107), 
         .D(n29182), .Z(clk_enable_400)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_520.init = 16'h55d5;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_521 (.A(resetn_c), .B(n13074), .C(n29124), 
         .D(n29127), .Z(clk_enable_402)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_521.init = 16'h5d55;
    LUT4 i2_3_lut_4_lut_4_lut_adj_522 (.A(resetn_c), .B(quad_set_complete_adj_149), 
         .C(n29134), .D(n29127), .Z(clk_enable_503)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i2_3_lut_4_lut_4_lut_adj_522.init = 16'hfddd;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_523 (.A(resetn_c), .B(n29213), .C(n29124), 
         .D(n29127), .Z(clk_enable_30)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // c:/s_links/sources/status_led.v(41[6:13])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_523.init = 16'h5d55;
    LUT4 i1_2_lut_rep_512 (.A(n2724), .B(spi_cmd_start_reg_N_746), .Z(n29240)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_2_lut_rep_512.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(n2724), .B(spi_cmd_start_reg_N_746), .C(n2713[4]), 
         .Z(n4606)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_513 (.A(n2713[7]), .B(n2713[3]), .Z(n29241)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_2_lut_rep_513.init = 16'heeee;
    LUT4 i1_3_lut_4_lut (.A(n2713[7]), .B(n2713[3]), .C(n2720), .D(n29318), 
         .Z(n5876)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_3_lut_4_lut.init = 16'hfe00;
    LUT4 i20046_3_lut_4_lut (.A(spi_byte_cnt[1]), .B(spi_byte_cnt[0]), .C(spi_byte_cnt[2]), 
         .D(spi_byte_cnt[3]), .Z(n21[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/s_links/sources/spi_ctrl.v(383[46:62])
    defparam i20046_3_lut_4_lut.init = 16'h7f80;
    LUT4 i20039_2_lut_3_lut (.A(spi_byte_cnt[1]), .B(spi_byte_cnt[0]), .C(spi_byte_cnt[2]), 
         .Z(n21[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(383[46:62])
    defparam i20039_2_lut_3_lut.init = 16'h7878;
    LUT4 i1_2_lut_rep_520 (.A(n2713[10]), .B(\address_7__N_549[1] ), .Z(n29248)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_520.init = 16'h8888;
    LUT4 i5936_3_lut_3_lut_3_lut (.A(n2713[10]), .B(\address_7__N_549[1] ), 
         .C(spi_cmd[15]), .Z(n10729)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B))) */ ;
    defparam i5936_3_lut_3_lut_3_lut.init = 16'h4c4c;
    FD1P3IX spi_byte_cnt_2505__i0 (.D(n21[0]), .SP(clk_enable_516), .CD(n29176), 
            .CK(clk), .Q(spi_byte_cnt[0]));   // c:/s_links/sources/spi_ctrl.v(383[46:62])
    defparam spi_byte_cnt_2505__i0.GSR = "ENABLED";
    LUT4 i5140_4_lut_4_lut (.A(n2713[10]), .B(\address_7__N_549[1] ), .C(n29073), 
         .D(spi_cmd[15]), .Z(address_7__N_359[0])) /* synthesis lut_function=(A ((D)+!B)+!A !(B (C))) */ ;
    defparam i5140_4_lut_4_lut.init = 16'hbf37;
    LUT4 i2215_3_lut_rep_524 (.A(spi_cmd_start_reg_N_745), .B(\address_7__N_549[1] ), 
         .C(n2713[10]), .Z(n29252)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i2215_3_lut_rep_524.init = 16'hcaca;
    FD1S3IX mem_rdata_update_206 (.D(n9633), .CK(clk), .CD(wr_en_N_355), 
            .Q(mem_rdata_update)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(79[9] 86[5])
    defparam mem_rdata_update_206.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_452_4_lut (.A(spi_cmd_start_reg_N_745), .B(\address_7__N_549[1] ), 
         .C(n2713[10]), .D(spi_cmd[15]), .Z(n29180)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_2_lut_rep_452_4_lut.init = 16'h00ca;
    LUT4 i60_4_lut_4_lut (.A(n29186), .B(n29269), .C(n2713[10]), .D(n26_adj_6703), 
         .Z(n38_adj_6704)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/s_links/sources/spi_ctrl.v(70[16:29])
    defparam i60_4_lut_4_lut.init = 16'h4f40;
    FD1P3IX mem_burst_cnt_2507__i0 (.D(n37[0]), .SP(clk_enable_309), .CD(n29179), 
            .CK(clk), .Q(mem_burst_cnt[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_2507__i0.GSR = "ENABLED";
    LUT4 i5179_4_lut_4_lut (.A(n29186), .B(clk_enable_366), .C(mem_rdata_update_N_729), 
         .D(\address_7__N_549[1] ), .Z(n9972)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B+!((D)+!C)))) */ ;   // c:/s_links/sources/spi_ctrl.v(70[16:29])
    defparam i5179_4_lut_4_lut.init = 16'h44f4;
    LUT4 i1_3_lut_rep_413 (.A(spi_addr[3]), .B(n27465), .C(n26928), .Z(n29141)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_3_lut_rep_413.init = 16'hfefe;
    LUT4 i1_2_lut_rep_398_4_lut (.A(spi_addr[3]), .B(n27465), .C(n26928), 
         .D(spi_cmd[1]), .Z(n29126)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i1_2_lut_rep_398_4_lut.init = 16'hfeff;
    LUT4 i14386_3_lut_4_lut (.A(wb_dat_o[3]), .B(n29186), .C(wb_dat_o[4]), 
         .D(\address_7__N_549[1] ), .Z(n19324)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i14386_3_lut_4_lut.init = 16'hfe00;
    LUT4 i22431_2_lut_3_lut_4_lut (.A(wb_dat_o[4]), .B(n29186), .C(\address_7__N_549[1] ), 
         .D(wb_dat_o[3]), .Z(n27601)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(255[32] 262[30])
    defparam i22431_2_lut_3_lut_4_lut.init = 16'hf0e0;
    PFUMX i23062 (.BLUT(n28765), .ALUT(n28764), .C0(spi_cmd_start_reg), 
          .Z(n28766));
    FD1P3AX mem_addr_2509__i0 (.D(n47[0]), .SP(clk_enable_516), .CK(clk), 
            .Q(spi_addr[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509__i0.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_534 (.A(spi_cmd[10]), .B(spi_cmd[12]), .C(spi_cmd[8]), 
         .Z(n29262)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_534.init = 16'hfefe;
    LUT4 i22448_2_lut_4_lut (.A(spi_cmd[10]), .B(spi_cmd[12]), .C(spi_cmd[8]), 
         .D(n22_adj_6705), .Z(n27618)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i22448_2_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(mem_burst_cnt[4]), .B(mem_burst_cnt[1]), .Z(n8)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(355[47:82])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i8772_3_lut_rep_345 (.A(n5874), .B(spi_addr_valid_N_732), .C(n5880), 
         .Z(n29073)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i8772_3_lut_rep_345.init = 16'hcece;
    PFUMX i5937 (.BLUT(n6901[1]), .ALUT(n10729), .C0(n27679), .Z(address_7__N_359[1]));
    LUT4 spi_xfer_done_I_10_2_lut_rep_538 (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .Z(n29266)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam spi_xfer_done_I_10_2_lut_rep_538.init = 16'h4444;
    LUT4 i15_1_lut_rep_408_2_lut_3_lut (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(spi_idle), .Z(n29136)) /* synthesis lut_function=(!(A (C)+!A (B+(C)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam i15_1_lut_rep_408_2_lut_3_lut.init = 16'h0b0b;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(n29318), .D(spi_idle), .Z(n4_adj_6706)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B+((D)+!C)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'h00b0;
    LUT4 spi_xfer_done_I_0_240_2_lut_rep_458_3_lut (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(spi_idle), .Z(n29186)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam spi_xfer_done_I_0_240_2_lut_rep_458_3_lut.init = 16'hf4f4;
    LUT4 wb_xfer_done_I_0_239_2_lut_3_lut_4_lut (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(\address_7__N_549[1] ), .D(spi_idle), .Z(wr_en_N_703)) /* synthesis lut_function=(A (C (D))+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam wb_xfer_done_I_0_239_2_lut_3_lut_4_lut.init = 16'hf040;
    LUT4 i1213_2_lut_rep_415_3_lut_4_lut (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(wb_dat_o[4]), .D(spi_idle), .Z(n29143)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam i1213_2_lut_rep_415_3_lut_4_lut.init = 16'hfff4;
    LUT4 i1_2_lut_rep_414_3_lut_4_lut (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(wb_dat_o[3]), .D(spi_idle), .Z(n29142)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam i1_2_lut_rep_414_3_lut_4_lut.init = 16'hfff4;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_adj_524 (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(n2724), .D(spi_idle), .Z(n27180)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B+((D)+!C)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam i1_2_lut_2_lut_3_lut_4_lut_adj_524.init = 16'h00b0;
    LUT4 i22413_2_lut_3_lut_4_lut (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(n29319), .D(spi_idle), .Z(n27578)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:62])
    defparam i22413_2_lut_3_lut_4_lut.init = 16'hfff4;
    LUT4 spi_cmd_start_I_15_2_lut_3_lut (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .C(spi_cmd_start_reg), .Z(spi_cmd_start)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(123[28:62])
    defparam spi_cmd_start_I_15_2_lut_3_lut.init = 16'hf2f2;
    LUT4 i22889_2_lut_rep_540 (.A(rd_en), .B(wr_en), .Z(n29268)) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i22889_2_lut_rep_540.init = 16'h1111;
    LUT4 n18805_bdd_3_lut_4_lut (.A(rd_en), .B(wr_en), .C(wb_sm), .D(\address_7__N_549[1] ), 
         .Z(n28767)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam n18805_bdd_3_lut_4_lut.init = 16'h0efe;
    LUT4 i1_2_lut_3_lut_adj_525 (.A(rd_en), .B(wr_en), .C(wb_sm), .Z(wb_cyc_i_N_339)) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_2_lut_3_lut_adj_525.init = 16'h0e0e;
    LUT4 i5003_2_lut_rep_541 (.A(spi_cmd[15]), .B(\address_7__N_549[1] ), 
         .Z(n29269)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/s_links/sources/spi_ctrl.v(307[24] 343[27])
    defparam i5003_2_lut_rep_541.init = 16'h4444;
    LUT4 i22873_2_lut_rep_459_3_lut (.A(spi_cmd[15]), .B(\address_7__N_549[1] ), 
         .C(n2713[10]), .Z(n29187)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(307[24] 343[27])
    defparam i22873_2_lut_rep_459_3_lut.init = 16'hbfbf;
    LUT4 i11_3_lut_4_lut (.A(spi_cmd[15]), .B(\address_7__N_549[1] ), .C(n2713[10]), 
         .D(n29308), .Z(clk_enable_504)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/s_links/sources/spi_ctrl.v(307[24] 343[27])
    defparam i11_3_lut_4_lut.init = 16'h4f40;
    LUT4 i22541_3_lut_4_lut (.A(\address_7__N_565[1] ), .B(n5874), .C(n5880), 
         .D(n5876), .Z(n6901[1])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i22541_3_lut_4_lut.init = 16'hf202;
    LUT4 i22460_2_lut_3_lut (.A(spi_addr_valid_N_732), .B(n29238), .C(n2720), 
         .Z(n27630)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i22460_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_adj_526 (.A(spi_cmd[15]), .B(n29252), .C(spi_data_valid_N_737), 
         .Z(clk_enable_474)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_3_lut_adj_526.init = 16'h4040;
    LUT4 i1_2_lut_adj_527 (.A(spi_byte_cnt[1]), .B(n26945), .Z(clk_enable_482)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_527.init = 16'h8888;
    LUT4 i2_4_lut (.A(spi_byte_cnt[2]), .B(n29180), .C(spi_byte_cnt[3]), 
         .D(spi_byte_cnt[0]), .Z(n26945)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i2_4_lut.init = 16'h0400;
    LUT4 i5_3_lut (.A(spi_byte_cnt[3]), .B(n10), .C(n29252), .Z(clk_enable_490)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i5_3_lut.init = 16'h4040;
    LUT4 i4_4_lut (.A(spi_cmd[15]), .B(spi_byte_cnt[1]), .C(spi_byte_cnt[0]), 
         .D(spi_byte_cnt[2]), .Z(n10)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i4_4_lut.init = 16'h0004;
    LUT4 i1_2_lut_adj_528 (.A(spi_byte_cnt[1]), .B(n26945), .Z(clk_enable_498)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_528.init = 16'h4444;
    LUT4 spi_xfer_done_N_706_bdd_3_lut_23041_4_lut (.A(n29266), .B(spi_idle), 
         .C(\address_7__N_549[1] ), .D(spi_cmd[15]), .Z(n28722)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:73])
    defparam spi_xfer_done_N_706_bdd_3_lut_23041_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_400_3_lut_4_lut (.A(n29266), .B(spi_idle), .C(wb_dat_o[3]), 
         .D(wb_dat_o[4]), .Z(n29128)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:73])
    defparam i1_2_lut_rep_400_3_lut_4_lut.init = 16'hfffe;
    LUT4 i14351_2_lut_rep_397_3_lut_4_lut (.A(n29266), .B(spi_idle), .C(\address_7__N_549[1] ), 
         .D(wb_dat_o[3]), .Z(n29125)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:73])
    defparam i14351_2_lut_rep_397_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i13996_3_lut_3_lut_4_lut (.A(n29266), .B(spi_idle), .C(\address_7__N_549[1] ), 
         .D(wb_dat_o[3]), .Z(rd_en_N_717)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:73])
    defparam i13996_3_lut_3_lut_4_lut.init = 16'hf010;
    LUT4 i2_3_lut_3_lut_3_lut_4_lut (.A(n29266), .B(spi_idle), .C(n4_adj_6707), 
         .D(n29187), .Z(n25453)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(135[28:73])
    defparam i2_3_lut_3_lut_3_lut_4_lut.init = 16'hf0f1;
    PFUMX i57 (.BLUT(n38_adj_6704), .ALUT(n32_adj_6708), .C0(n27675), 
          .Z(rd_en_N_710));
    LUT4 i1261_2_lut_rep_551 (.A(\address_7__N_549[1] ), .B(n2713[4]), .Z(n29279)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1261_2_lut_rep_551.init = 16'h8888;
    LUT4 i5259_2_lut_3_lut (.A(\address_7__N_549[1] ), .B(n2713[4]), .C(spi_cmd_cnt), 
         .Z(clk_enable_525)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i5259_2_lut_3_lut.init = 16'h8080;
    LUT4 i22962_2_lut_4_lut (.A(n5874), .B(spi_addr_valid_N_732), .C(n5880), 
         .D(n29248), .Z(n27679)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B+(D))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i22962_2_lut_4_lut.init = 16'hffce;
    LUT4 i22935_2_lut_3_lut (.A(\address_7__N_549[1] ), .B(n2713[4]), .C(spi_cmd_cnt), 
         .Z(clk_enable_279)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i22935_2_lut_3_lut.init = 16'h0808;
    LUT4 mem_addr_2509_mux_6_i2_3_lut (.A(wb_dat_o[1]), .B(n37_adj_6725[1]), 
         .C(n7083), .Z(n47[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509_mux_6_i2_3_lut.init = 16'hcaca;
    LUT4 i3_3_lut_4_lut (.A(spi_cmd[15]), .B(n29319), .C(n2713[10]), .D(n2713[4]), 
         .Z(n8_adj_6709)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i3_3_lut_4_lut.init = 16'h0008;
    LUT4 i13721_2_lut (.A(mem_rdata[0]), .B(mem_wr_N_726), .Z(n672[0])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(358[46:63])
    defparam i13721_2_lut.init = 16'hbbbb;
    LUT4 mem_addr_2509_mux_6_i3_3_lut (.A(wb_dat_o[2]), .B(n37_adj_6725[2]), 
         .C(n7083), .Z(n47[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509_mux_6_i3_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut (.A(n19198), .B(n26923), .C(mem_burst_cnt[4]), .D(mem_burst_cnt[1]), 
         .Z(mem_wr_N_726)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/s_links/sources/spi_ctrl.v(355[47:82])
    defparam i3_4_lut.init = 16'hfffd;
    LUT4 mem_addr_2509_mux_6_i4_3_lut (.A(wb_dat_o[3]), .B(n37_adj_6725[3]), 
         .C(n7083), .Z(n47[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509_mux_6_i4_3_lut.init = 16'hcaca;
    LUT4 mem_addr_2509_mux_6_i5_3_lut (.A(wb_dat_o[4]), .B(n37_adj_6725[4]), 
         .C(n7083), .Z(n47[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509_mux_6_i5_3_lut.init = 16'hcaca;
    LUT4 mem_addr_2509_mux_6_i6_3_lut (.A(wb_dat_o[5]), .B(n37_adj_6725[5]), 
         .C(n7083), .Z(n47[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509_mux_6_i6_3_lut.init = 16'hcaca;
    LUT4 mem_addr_2509_mux_6_i7_3_lut (.A(wb_dat_o[6]), .B(n37_adj_6725[6]), 
         .C(n7083), .Z(n47[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509_mux_6_i7_3_lut.init = 16'hcaca;
    LUT4 i14271_2_lut (.A(mem_burst_cnt[0]), .B(mem_burst_cnt[2]), .Z(n19198)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14271_2_lut.init = 16'h8888;
    LUT4 mem_addr_2509_mux_6_i8_3_lut (.A(wb_dat_o[7]), .B(n37_adj_6725[7]), 
         .C(n7083), .Z(n47[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509_mux_6_i8_3_lut.init = 16'hcaca;
    CCU2D mem_burst_cnt_2507_add_4_9 (.A0(mem_burst_cnt[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25199), .S0(n37[7]));   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_2507_add_4_9.INIT0 = 16'hfaaa;
    defparam mem_burst_cnt_2507_add_4_9.INIT1 = 16'h0000;
    defparam mem_burst_cnt_2507_add_4_9.INJECT1_0 = "NO";
    defparam mem_burst_cnt_2507_add_4_9.INJECT1_1 = "NO";
    CCU2D mem_burst_cnt_2507_add_4_7 (.A0(mem_burst_cnt[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(mem_burst_cnt[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n25198), .COUT(n25199), .S0(n37[5]), 
          .S1(n37[6]));   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_2507_add_4_7.INIT0 = 16'hfaaa;
    defparam mem_burst_cnt_2507_add_4_7.INIT1 = 16'hfaaa;
    defparam mem_burst_cnt_2507_add_4_7.INJECT1_0 = "NO";
    defparam mem_burst_cnt_2507_add_4_7.INJECT1_1 = "NO";
    CCU2D mem_burst_cnt_2507_add_4_5 (.A0(mem_burst_cnt[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(mem_burst_cnt[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n25197), .COUT(n25198), .S0(n37[3]), 
          .S1(n37[4]));   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_2507_add_4_5.INIT0 = 16'hfaaa;
    defparam mem_burst_cnt_2507_add_4_5.INIT1 = 16'hfaaa;
    defparam mem_burst_cnt_2507_add_4_5.INJECT1_0 = "NO";
    defparam mem_burst_cnt_2507_add_4_5.INJECT1_1 = "NO";
    CCU2D mem_burst_cnt_2507_add_4_3 (.A0(mem_burst_cnt[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(mem_burst_cnt[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n25196), .COUT(n25197), .S0(n37[1]), 
          .S1(n37[2]));   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_2507_add_4_3.INIT0 = 16'hfaaa;
    defparam mem_burst_cnt_2507_add_4_3.INIT1 = 16'hfaaa;
    defparam mem_burst_cnt_2507_add_4_3.INJECT1_0 = "NO";
    defparam mem_burst_cnt_2507_add_4_3.INJECT1_1 = "NO";
    CCU2D mem_burst_cnt_2507_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(mem_burst_cnt[0]), .B1(n19198), .C1(n8), 
          .D1(n26923), .COUT(n25196), .S1(n37[0]));   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_2507_add_4_1.INIT0 = 16'hF000;
    defparam mem_burst_cnt_2507_add_4_1.INIT1 = 16'h5559;
    defparam mem_burst_cnt_2507_add_4_1.INJECT1_0 = "NO";
    defparam mem_burst_cnt_2507_add_4_1.INJECT1_1 = "NO";
    CCU2D mem_addr_2509_add_4_9 (.A0(spi_addr[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25195), .S0(n37_adj_6725[7]));   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509_add_4_9.INIT0 = 16'hfaaa;
    defparam mem_addr_2509_add_4_9.INIT1 = 16'h0000;
    defparam mem_addr_2509_add_4_9.INJECT1_0 = "NO";
    defparam mem_addr_2509_add_4_9.INJECT1_1 = "NO";
    CCU2D mem_addr_2509_add_4_7 (.A0(spi_addr[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_addr[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25194), .COUT(n25195), .S0(n37_adj_6725[5]), 
          .S1(n37_adj_6725[6]));   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509_add_4_7.INIT0 = 16'hfaaa;
    defparam mem_addr_2509_add_4_7.INIT1 = 16'hfaaa;
    defparam mem_addr_2509_add_4_7.INJECT1_0 = "NO";
    defparam mem_addr_2509_add_4_7.INJECT1_1 = "NO";
    CCU2D mem_addr_2509_add_4_5 (.A0(spi_addr[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_addr[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25193), .COUT(n25194), .S0(n37_adj_6725[3]), 
          .S1(n37_adj_6725[4]));   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509_add_4_5.INIT0 = 16'hfaaa;
    defparam mem_addr_2509_add_4_5.INIT1 = 16'hfaaa;
    defparam mem_addr_2509_add_4_5.INJECT1_0 = "NO";
    defparam mem_addr_2509_add_4_5.INJECT1_1 = "NO";
    LUT4 i3_4_lut_adj_529 (.A(mem_burst_cnt[6]), .B(mem_burst_cnt[5]), .C(mem_burst_cnt[3]), 
         .D(mem_burst_cnt[7]), .Z(n26923)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(355[47:82])
    defparam i3_4_lut_adj_529.init = 16'hfffe;
    CCU2D mem_addr_2509_add_4_3 (.A0(spi_addr[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_addr[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n25192), .COUT(n25193), .S0(n37_adj_6725[1]), 
          .S1(n37_adj_6725[2]));   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509_add_4_3.INIT0 = 16'hfaaa;
    defparam mem_addr_2509_add_4_3.INIT1 = 16'hfaaa;
    defparam mem_addr_2509_add_4_3.INJECT1_0 = "NO";
    defparam mem_addr_2509_add_4_3.INJECT1_1 = "NO";
    CCU2D mem_addr_2509_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(spi_addr[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n25192), .S1(n37_adj_6725[0]));   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509_add_4_1.INIT0 = 16'hF000;
    defparam mem_addr_2509_add_4_1.INIT1 = 16'h0555;
    defparam mem_addr_2509_add_4_1.INJECT1_0 = "NO";
    defparam mem_addr_2509_add_4_1.INJECT1_1 = "NO";
    LUT4 i14021_2_lut_3_lut (.A(spi_cmd_start_reg_N_745), .B(n2724), .C(n2713[4]), 
         .Z(n18948)) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;
    defparam i14021_2_lut_3_lut.init = 16'h0e0e;
    LUT4 i11_3_lut_4_lut_adj_530 (.A(spi_cmd_start_reg_N_745), .B(n2724), 
         .C(n2713[4]), .D(\address_7__N_549[1] ), .Z(clk_enable_507)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam i11_3_lut_4_lut_adj_530.init = 16'hfe0e;
    FD1P3AX spi_cmd_i0_i15 (.D(wb_dat_o[7]), .SP(clk_enable_279), .CK(clk), 
            .Q(spi_cmd[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i15.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i14 (.D(wb_dat_o[6]), .SP(clk_enable_279), .CK(clk), 
            .Q(spi_cmd[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i14.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i13 (.D(wb_dat_o[5]), .SP(clk_enable_279), .CK(clk), 
            .Q(spi_cmd[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i13.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i12 (.D(wb_dat_o[4]), .SP(clk_enable_279), .CK(clk), 
            .Q(spi_cmd[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i12.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i11 (.D(wb_dat_o[3]), .SP(clk_enable_279), .CK(clk), 
            .Q(spi_cmd[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i11.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i10 (.D(wb_dat_o[2]), .SP(clk_enable_279), .CK(clk), 
            .Q(spi_cmd[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i10.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i9 (.D(wb_dat_o[1]), .SP(clk_enable_279), .CK(clk), 
            .Q(spi_cmd[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i9.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i8 (.D(wb_dat_o[0]), .SP(clk_enable_279), .CK(clk), 
            .Q(spi_cmd[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i8.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i7 (.D(wb_dat_o[7]), .SP(clk_enable_525), .CK(clk), 
            .Q(spi_cmd[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i7.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i6 (.D(wb_dat_o[6]), .SP(clk_enable_525), .CK(clk), 
            .Q(spi_cmd[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i6.GSR = "ENABLED";
    PFUMX i59 (.BLUT(n36), .ALUT(rd_en_N_717), .C0(n2720), .Z(n26_adj_6703));
    FD1P3AX spi_cmd_i0_i5 (.D(wb_dat_o[5]), .SP(clk_enable_525), .CK(clk), 
            .Q(spi_cmd[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i5.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i4 (.D(wb_dat_o[4]), .SP(clk_enable_525), .CK(clk), 
            .Q(spi_cmd[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i4.GSR = "ENABLED";
    FD1P3AY spi_cmd_i0_i3 (.D(wb_dat_o[3]), .SP(clk_enable_525), .CK(clk), 
            .Q(spi_cmd[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i3.GSR = "ENABLED";
    FD1P3AX spi_cmd_i0_i2 (.D(wb_dat_o[2]), .SP(clk_enable_525), .CK(clk), 
            .Q(spi_cmd[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i2.GSR = "ENABLED";
    PFUMX i23039 (.BLUT(n29136), .ALUT(n28722), .C0(wb_dat_o[4]), .Z(n28723));
    LUT4 i20032_2_lut (.A(spi_byte_cnt[1]), .B(spi_byte_cnt[0]), .Z(n21[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/spi_ctrl.v(383[46:62])
    defparam i20032_2_lut.init = 16'h6666;
    LUT4 i4779_3_lut_4_lut (.A(resetn_c), .B(n29114), .C(n29213), .D(reset_r_N_4474), 
         .Z(clk_enable_20)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(D))) */ ;
    defparam i4779_3_lut_4_lut.init = 16'h7f00;
    FD1P3AY spi_cmd_i0_i1 (.D(wb_dat_o[1]), .SP(clk_enable_525), .CK(clk), 
            .Q(spi_cmd[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i1.GSR = "ENABLED";
    FD1P3AY spi_cmd_i0_i0 (.D(wb_dat_o[0]), .SP(clk_enable_525), .CK(clk), 
            .Q(spi_cmd[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i0.GSR = "ENABLED";
    FD1P3IX mem_burst_cnt_2507__i2 (.D(n37[2]), .SP(clk_enable_309), .CD(n29179), 
            .CK(clk), .Q(mem_burst_cnt[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_2507__i2.GSR = "ENABLED";
    FD1P3IX mem_burst_cnt_2507__i1 (.D(n37[1]), .SP(clk_enable_309), .CD(n29179), 
            .CK(clk), .Q(mem_burst_cnt[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(385[50:67])
    defparam mem_burst_cnt_2507__i1.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(spi_cmd_start_reg_N_745), .B(n29186), .C(\address_7__N_565[1] ), 
         .D(n18), .Z(n26429)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut.init = 16'hce0a;
    LUT4 i2_4_lut_adj_531 (.A(\address_7__N_549[1] ), .B(n2724), .C(n15), 
         .D(n29187), .Z(n18)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+!(D))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i2_4_lut_adj_531.init = 16'hecff;
    LUT4 i1_4_lut_adj_532 (.A(n29318), .B(n2713[11]), .C(n13622), .D(n2713[7]), 
         .Z(n15)) /* synthesis lut_function=(A (B+(D))+!A (B+(C+(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_532.init = 16'hffdc;
    LUT4 i1_4_lut_adj_533 (.A(spi_cmd_start), .B(n29268), .C(\address_7__N_549[1] ), 
         .D(wb_sm), .Z(n30)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_533.init = 16'ha088;
    LUT4 i4_2_lut (.A(n2713[3]), .B(n2720), .Z(n13622)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i4_2_lut.init = 16'heeee;
    FD1P3AX wr_data_i0_i1 (.D(n672[1]), .SP(clk_enable_366), .CK(clk), 
            .Q(wr_data[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i1.GSR = "ENABLED";
    FD1P3AX wr_data_i0_i2 (.D(n672[2]), .SP(clk_enable_366), .CK(clk), 
            .Q(wr_data[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i2.GSR = "ENABLED";
    FD1P3AX wr_data_i0_i3 (.D(n672[3]), .SP(clk_enable_366), .CK(clk), 
            .Q(wr_data[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i3.GSR = "ENABLED";
    FD1P3AX wr_data_i0_i4 (.D(n672[4]), .SP(clk_enable_366), .CK(clk), 
            .Q(wr_data[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i4.GSR = "ENABLED";
    FD1P3AX wr_data_i0_i5 (.D(n672[5]), .SP(clk_enable_366), .CK(clk), 
            .Q(wr_data[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i5.GSR = "ENABLED";
    FD1P3AX wr_data_i0_i6 (.D(n672[6]), .SP(clk_enable_366), .CK(clk), 
            .Q(wr_data[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i6.GSR = "ENABLED";
    FD1P3AX wr_data_i0_i7 (.D(n672[7]), .SP(clk_enable_366), .CK(clk), 
            .Q(wr_data[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam wr_data_i0_i7.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i2 (.D(n9429), .CK(clk), .Q(spi_cmd_start_reg_N_746));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i2.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i3 (.D(n26319), .CK(clk), .Q(n2713[2]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i3.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i4 (.D(n9988), .CK(clk), .Q(n2713[3]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i4.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i5 (.D(n9986), .CK(clk), .Q(n2713[4]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i5.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i6 (.D(n29279), .CK(clk), .Q(n2724));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i6.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i7 (.D(n25364), .CK(clk), .Q(n2713[6]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i7.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i8 (.D(n9982), .CK(clk), .Q(n2713[7]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i8.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i9 (.D(n9980), .CK(clk), .Q(spi_addr_valid_N_732));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i9.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i10 (.D(n25453), .CK(clk), .Q(n2720));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i10.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i11 (.D(n9976), .CK(clk), .Q(n2713[10]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i11.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i12 (.D(n13_adj_6718), .CK(clk), .Q(n2713[11]));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i12.GSR = "ENABLED";
    FD1S3AX main_sm_FSM_i13 (.D(n9972), .CK(clk), .Q(mem_rdata_update_N_729));   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam main_sm_FSM_i13.GSR = "ENABLED";
    FD1P3IX spi_data__i1 (.D(wb_dat_o[1]), .SP(clk_enable_474), .CD(n7710), 
            .CK(clk), .Q(\spi_data[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i1.GSR = "ENABLED";
    FD1P3IX spi_data__i2 (.D(wb_dat_o[2]), .SP(clk_enable_474), .CD(n7710), 
            .CK(clk), .Q(\spi_data[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i2.GSR = "ENABLED";
    FD1P3IX spi_data__i3 (.D(wb_dat_o[3]), .SP(clk_enable_474), .CD(n7710), 
            .CK(clk), .Q(\spi_data[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i3.GSR = "ENABLED";
    FD1P3IX spi_data__i4 (.D(wb_dat_o[4]), .SP(clk_enable_474), .CD(n7710), 
            .CK(clk), .Q(\spi_data[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i4.GSR = "ENABLED";
    FD1P3IX spi_data__i5 (.D(wb_dat_o[5]), .SP(clk_enable_474), .CD(n7710), 
            .CK(clk), .Q(\spi_data[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i5.GSR = "ENABLED";
    FD1P3IX spi_data__i6 (.D(wb_dat_o[6]), .SP(clk_enable_474), .CD(n7710), 
            .CK(clk), .Q(\spi_data[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i6.GSR = "ENABLED";
    FD1P3IX spi_data__i7 (.D(wb_dat_o[7]), .SP(clk_enable_474), .CD(n7710), 
            .CK(clk), .Q(\spi_data[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i7.GSR = "ENABLED";
    FD1P3IX spi_data__i8 (.D(wb_dat_o[0]), .SP(clk_enable_482), .CD(n7710), 
            .CK(clk), .Q(\spi_data[8] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i8.GSR = "ENABLED";
    FD1P3IX spi_data__i9 (.D(wb_dat_o[1]), .SP(clk_enable_482), .CD(n7710), 
            .CK(clk), .Q(\spi_data[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i9.GSR = "ENABLED";
    FD1P3IX spi_data__i10 (.D(wb_dat_o[2]), .SP(clk_enable_482), .CD(n7710), 
            .CK(clk), .Q(\spi_data[10] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i10.GSR = "ENABLED";
    FD1P3IX spi_data__i11 (.D(wb_dat_o[3]), .SP(clk_enable_482), .CD(n7710), 
            .CK(clk), .Q(\spi_data[11] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i11.GSR = "ENABLED";
    FD1P3IX spi_data__i12 (.D(wb_dat_o[4]), .SP(clk_enable_482), .CD(n7710), 
            .CK(clk), .Q(\spi_data[12] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i12.GSR = "ENABLED";
    FD1P3IX spi_data__i13 (.D(wb_dat_o[5]), .SP(clk_enable_482), .CD(n7710), 
            .CK(clk), .Q(\spi_data[13] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i13.GSR = "ENABLED";
    FD1P3IX spi_data__i14 (.D(wb_dat_o[6]), .SP(clk_enable_482), .CD(n7710), 
            .CK(clk), .Q(\spi_data[14] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i14.GSR = "ENABLED";
    FD1P3IX spi_data__i15 (.D(wb_dat_o[7]), .SP(clk_enable_482), .CD(n7710), 
            .CK(clk), .Q(\spi_data[15] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i15.GSR = "ENABLED";
    FD1P3IX spi_data__i16 (.D(wb_dat_o[0]), .SP(clk_enable_490), .CD(n7710), 
            .CK(clk), .Q(\spi_data[16] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i16.GSR = "ENABLED";
    FD1P3IX spi_data__i17 (.D(wb_dat_o[1]), .SP(clk_enable_490), .CD(n7710), 
            .CK(clk), .Q(\spi_data[17] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i17.GSR = "ENABLED";
    FD1P3IX spi_data__i18 (.D(wb_dat_o[2]), .SP(clk_enable_490), .CD(n7710), 
            .CK(clk), .Q(\spi_data[18] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i18.GSR = "ENABLED";
    FD1P3IX spi_data__i19 (.D(wb_dat_o[3]), .SP(clk_enable_490), .CD(n7710), 
            .CK(clk), .Q(\spi_data[19] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i19.GSR = "ENABLED";
    FD1P3IX spi_data__i20 (.D(wb_dat_o[4]), .SP(clk_enable_490), .CD(n7710), 
            .CK(clk), .Q(\spi_data[20] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i20.GSR = "ENABLED";
    FD1P3IX spi_data__i21 (.D(wb_dat_o[5]), .SP(clk_enable_490), .CD(n7710), 
            .CK(clk), .Q(\spi_data[21] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i21.GSR = "ENABLED";
    FD1P3IX spi_data__i22 (.D(wb_dat_o[6]), .SP(clk_enable_490), .CD(n7710), 
            .CK(clk), .Q(\spi_data[22] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i22.GSR = "ENABLED";
    FD1P3IX spi_data__i23 (.D(wb_dat_o[7]), .SP(clk_enable_490), .CD(n7710), 
            .CK(clk), .Q(\spi_data[23] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i23.GSR = "ENABLED";
    FD1P3IX spi_data__i24 (.D(wb_dat_o[0]), .SP(clk_enable_498), .CD(n7710), 
            .CK(clk), .Q(\spi_data[24] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i24.GSR = "ENABLED";
    FD1P3IX spi_data__i25 (.D(wb_dat_o[1]), .SP(clk_enable_498), .CD(n7710), 
            .CK(clk), .Q(\spi_data[25] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i25.GSR = "ENABLED";
    FD1P3IX spi_data__i26 (.D(wb_dat_o[2]), .SP(clk_enable_498), .CD(n7710), 
            .CK(clk), .Q(\spi_data[26] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i26.GSR = "ENABLED";
    FD1P3IX spi_data__i27 (.D(wb_dat_o[3]), .SP(clk_enable_498), .CD(n7710), 
            .CK(clk), .Q(\spi_data[27] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i27.GSR = "ENABLED";
    FD1P3IX spi_data__i28 (.D(wb_dat_o[4]), .SP(clk_enable_498), .CD(n7710), 
            .CK(clk), .Q(\spi_data[28] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i28.GSR = "ENABLED";
    FD1P3IX spi_data__i29 (.D(wb_dat_o[5]), .SP(clk_enable_498), .CD(n7710), 
            .CK(clk), .Q(\spi_data[29] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i29.GSR = "ENABLED";
    FD1P3IX spi_data__i30 (.D(wb_dat_o[6]), .SP(clk_enable_498), .CD(n7710), 
            .CK(clk), .Q(\spi_data[30] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i30.GSR = "ENABLED";
    FD1P3IX spi_data__i31 (.D(wb_dat_o[7]), .SP(clk_enable_498), .CD(n7710), 
            .CK(clk), .Q(\spi_data[31] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data__i31.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_580 (.A(n2720), .B(spi_cmd_start_reg_N_745), .Z(n29308)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_2_lut_rep_580.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_534 (.A(n2720), .B(spi_cmd_start_reg_N_745), 
         .C(n2713[10]), .Z(n18908)) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_2_lut_3_lut_adj_534.init = 16'h0e0e;
    FD1S3AX address_i2 (.D(address_7__N_359[1]), .CK(clk), .Q(\address[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam address_i2.GSR = "ENABLED";
    FD1S3IX mem_wr_219 (.D(mem_wr_N_726), .CK(clk), .CD(n29187), .Q(mem_wr)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam mem_wr_219.GSR = "ENABLED";
    FD1P3IX spi_data_valid_226 (.D(spi_data_valid_N_737), .SP(clk_enable_504), 
            .CD(n18908), .CK(clk), .Q(spi_data_valid)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_data_valid_226.GSR = "ENABLED";
    FD1P3IX spi_cmd_valid_223 (.D(spi_cmd_cnt), .SP(clk_enable_507), .CD(n18948), 
            .CK(clk), .Q(spi_cmd_valid)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_valid_223.GSR = "ENABLED";
    LUT4 i3_4_lut_adj_535 (.A(spi_cmd[5]), .B(spi_cmd[9]), .C(spi_cmd[3]), 
         .D(spi_cmd[6]), .Z(n22_adj_6705)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_535.init = 16'hfffe;
    LUT4 i1_4_lut_adj_536 (.A(n4606), .B(n29173), .C(\address_7__N_549[1] ), 
         .D(n27578), .Z(n36)) /* synthesis lut_function=(!(A+!(B (C)+!B !((D)+!C)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_536.init = 16'h4050;
    LUT4 i3_4_lut_adj_537 (.A(spi_cmd[11]), .B(spi_cmd[7]), .C(spi_cmd[13]), 
         .D(spi_cmd[14]), .Z(n31_adj_150)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_537.init = 16'hfffe;
    LUT4 wb_xfer_done_I_0_242_2_lut_rep_590 (.A(\address_7__N_549[1] ), .B(wb_dat_o[3]), 
         .Z(n29318)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_ctrl.v(288[31:57])
    defparam wb_xfer_done_I_0_242_2_lut_rep_590.init = 16'h8888;
    LUT4 i5193_4_lut_4_lut (.A(\address_7__N_549[1] ), .B(wb_dat_o[3]), 
         .C(n2713[3]), .D(n2713[4]), .Z(n9986)) /* synthesis lut_function=(A (B (C))+!A (D)) */ ;   // c:/s_links/sources/spi_ctrl.v(288[31:57])
    defparam i5193_4_lut_4_lut.init = 16'hd580;
    LUT4 i792_2_lut_3_lut (.A(\address_7__N_549[1] ), .B(wb_dat_o[3]), .C(n2720), 
         .Z(n2775)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(288[31:57])
    defparam i792_2_lut_3_lut.init = 16'h8080;
    LUT4 spi_xfer_done_bdd_3_lut_3_lut (.A(\address_7__N_549[1] ), .B(wb_dat_o[3]), 
         .C(wb_dat_o[4]), .Z(n28855)) /* synthesis lut_function=(A (B+!(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(288[31:57])
    defparam spi_xfer_done_bdd_3_lut_3_lut.init = 16'h8a8a;
    LUT4 spi_xfer_done_bdd_2_lut_3_lut (.A(\address_7__N_549[1] ), .B(wb_dat_o[3]), 
         .C(n2713[7]), .Z(n28854)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(288[31:57])
    defparam spi_xfer_done_bdd_2_lut_3_lut.init = 16'h0808;
    LUT4 wb_xfer_done_I_0_238_2_lut_rep_591 (.A(\address_7__N_549[1] ), .B(wb_dat_o[4]), 
         .Z(n29319)) /* synthesis lut_function=(A (B)) */ ;   // c:/s_links/sources/spi_ctrl.v(347[31:57])
    defparam wb_xfer_done_I_0_238_2_lut_rep_591.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_538 (.A(\address_7__N_549[1] ), .B(wb_dat_o[4]), 
         .C(n2713[11]), .Z(n6_adj_6720)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(347[31:57])
    defparam i1_2_lut_3_lut_adj_538.init = 16'h7070;
    LUT4 i1_2_lut_rep_388_3_lut_4_lut_4_lut (.A(\address_7__N_549[1] ), .B(wb_dat_o[4]), 
         .C(n29186), .D(wb_dat_o[3]), .Z(n29116)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(347[31:57])
    defparam i1_2_lut_rep_388_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\address_7__N_549[1] ), .B(wb_dat_o[4]), 
         .C(n2713[11]), .D(spi_cmd[15]), .Z(clk_enable_366)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(347[31:57])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i58_3_lut (.A(n28856), .B(n30), .C(spi_cmd_start_reg_N_745), 
         .Z(n32_adj_6708)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i58_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_539 (.A(spi_cmd_start_reg_N_745), .B(n2713[10]), .Z(n7710)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_adj_539.init = 16'h2222;
    LUT4 i22802_4_lut (.A(spi_byte_cnt[1]), .B(spi_byte_cnt[2]), .C(spi_byte_cnt[3]), 
         .D(spi_byte_cnt[0]), .Z(spi_data_valid_N_737)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/s_links/sources/spi_ctrl.v(331[12:16])
    defparam i22802_4_lut.init = 16'h0004;
    LUT4 i2_3_lut_4_lut (.A(n29319), .B(n29125), .C(n4_adj_6721), .D(n2713[7]), 
         .Z(n25364)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i2_3_lut_4_lut.init = 16'hf2f0;
    LUT4 i1_2_lut_adj_540 (.A(wr_en), .B(wb_sm), .Z(wb_we_i_N_344)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam i1_2_lut_adj_540.init = 16'h2222;
    LUT4 i20030_1_lut (.A(spi_byte_cnt[0]), .Z(n21[0])) /* synthesis lut_function=(!(A)) */ ;   // c:/s_links/sources/spi_ctrl.v(383[46:62])
    defparam i20030_1_lut.init = 16'h5555;
    LUT4 i22963_4_lut (.A(spi_cmd_start_reg_N_745), .B(n2713[10]), .C(n2720), 
         .D(n29241), .Z(n27675)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i22963_4_lut.init = 16'habaa;
    LUT4 i13656_2_lut (.A(mem_rdata[1]), .B(mem_wr_N_726), .Z(n672[1])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(358[46:63])
    defparam i13656_2_lut.init = 16'hbbbb;
    FD1P3AX mem_addr_2509__i1 (.D(n47[1]), .SP(clk_enable_516), .CK(clk), 
            .Q(spi_addr[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509__i1.GSR = "ENABLED";
    LUT4 i13655_2_lut (.A(mem_rdata[2]), .B(mem_wr_N_726), .Z(n672[2])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(358[46:63])
    defparam i13655_2_lut.init = 16'hbbbb;
    LUT4 i13654_2_lut (.A(mem_rdata[3]), .B(mem_wr_N_726), .Z(n672[3])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(358[46:63])
    defparam i13654_2_lut.init = 16'hbbbb;
    LUT4 i13653_2_lut (.A(mem_rdata[4]), .B(mem_wr_N_726), .Z(n672[4])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(358[46:63])
    defparam i13653_2_lut.init = 16'hbbbb;
    LUT4 i13646_2_lut (.A(mem_rdata[5]), .B(mem_wr_N_726), .Z(n672[5])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(358[46:63])
    defparam i13646_2_lut.init = 16'hbbbb;
    LUT4 i13645_2_lut (.A(mem_rdata[6]), .B(mem_wr_N_726), .Z(n672[6])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(358[46:63])
    defparam i13645_2_lut.init = 16'hbbbb;
    LUT4 i13644_2_lut (.A(mem_rdata[7]), .B(mem_wr_N_726), .Z(n672[7])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/spi_ctrl.v(358[46:63])
    defparam i13644_2_lut.init = 16'hbbbb;
    LUT4 i9241_3_lut (.A(spi_cmd_start_reg_N_745), .B(spi_idle_N_747), .C(spi_idle), 
         .Z(n14197)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(130[11] 133[31])
    defparam i9241_3_lut.init = 16'hdcdc;
    LUT4 i4662_4_lut (.A(spi_cmd_start_reg_N_746), .B(\address_7__N_565[1] ), 
         .C(\address_7__N_549[1] ), .D(spi_cmd_start_reg_N_745), .Z(n9429)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i4662_4_lut.init = 16'hce0a;
    LUT4 i2_4_lut_adj_541 (.A(n2713[2]), .B(n4_adj_6722), .C(spi_cmd_start_reg_N_746), 
         .D(\address_7__N_549[1] ), .Z(n26319)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i2_4_lut_adj_541.init = 16'hfcee;
    LUT4 i1_4_lut_adj_542 (.A(n2713[3]), .B(spi_cmd_cnt), .C(n29116), 
         .D(n27180), .Z(n4_adj_6722)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A !(B+!(D))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_542.init = 16'hb3a0;
    LUT4 i5195_4_lut (.A(n2713[3]), .B(\address_7__N_549[1] ), .C(n19324), 
         .D(n2713[2]), .Z(n9988)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i5195_4_lut.init = 16'hce0a;
    LUT4 i5_3_lut_adj_543 (.A(spi_cmd[4]), .B(n10_adj_6723), .C(spi_addr[5]), 
         .Z(n26928)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i5_3_lut_adj_543.init = 16'hfefe;
    LUT4 i1_4_lut_adj_544 (.A(spi_cmd_cnt), .B(n2713[6]), .C(n27180), 
         .D(\address_7__N_549[1] ), .Z(n4_adj_6721)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_544.init = 16'ha0ec;
    LUT4 i4_4_lut_adj_545 (.A(spi_addr[6]), .B(spi_addr[4]), .C(spi_cmd[15]), 
         .D(spi_addr[7]), .Z(n10_adj_6723)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i4_4_lut_adj_545.init = 16'hffef;
    LUT4 i5189_4_lut (.A(n2713[7]), .B(\address_7__N_549[1] ), .C(n19324), 
         .D(n2713[6]), .Z(n9982)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i5189_4_lut.init = 16'hce0a;
    LUT4 i5187_4_lut (.A(spi_addr_valid_N_732), .B(n2713[7]), .C(\address_7__N_549[1] ), 
         .D(n4_adj_6706), .Z(n9980)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i5187_4_lut.init = 16'hce0a;
    LUT4 i1_4_lut_adj_546 (.A(n29238), .B(n12), .C(n29241), .D(n27601), 
         .Z(n5874)) /* synthesis lut_function=(A+(B+!((D)+!C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_546.init = 16'heefe;
    LUT4 i1_4_lut_adj_547 (.A(wr_en_N_703), .B(n2720), .C(n6_adj_6720), 
         .D(n29318), .Z(n12)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C)))) */ ;
    defparam i1_4_lut_adj_547.init = 16'h5054;
    LUT4 i1_4_lut_adj_548 (.A(n29269), .B(n2720), .C(spi_addr_valid_N_732), 
         .D(n29125), .Z(n4_adj_6707)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((D)+!B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_548.init = 16'ha0ec;
    LUT4 i1_4_lut_adj_549 (.A(n4606), .B(n2713[10]), .C(n4_adj_6724), 
         .D(\address_7__N_549[1] ), .Z(n5880)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_549.init = 16'hfafe;
    LUT4 i2_3_lut (.A(n29262), .B(n31_adj_150), .C(n22_adj_6705), .Z(n27465)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam i2_3_lut.init = 16'hfefe;
    FD1P3AX mem_addr_2509__i2 (.D(n47[2]), .SP(clk_enable_516), .CK(clk), 
            .Q(spi_addr[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509__i2.GSR = "ENABLED";
    FD1P3AX mem_addr_2509__i3 (.D(n47[3]), .SP(clk_enable_516), .CK(clk), 
            .Q(spi_addr[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509__i3.GSR = "ENABLED";
    FD1P3AX mem_addr_2509__i4 (.D(n47[4]), .SP(clk_enable_516), .CK(clk), 
            .Q(spi_addr[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509__i4.GSR = "ENABLED";
    FD1P3AX mem_addr_2509__i5 (.D(n47[5]), .SP(clk_enable_516), .CK(clk), 
            .Q(spi_addr[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509__i5.GSR = "ENABLED";
    FD1P3AX mem_addr_2509__i6 (.D(n47[6]), .SP(clk_enable_516), .CK(clk), 
            .Q(spi_addr[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509__i6.GSR = "ENABLED";
    FD1P3AX mem_addr_2509__i7 (.D(n47[7]), .SP(clk_enable_516), .CK(clk), 
            .Q(spi_addr[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509__i7.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_550 (.A(\address_7__N_549[1] ), .B(n2713[11]), .C(n13568), 
         .D(n29143), .Z(n4_adj_6724)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_550.init = 16'ha8a0;
    LUT4 i3_4_lut_adj_551 (.A(n29128), .B(n29142), .C(n29241), .D(n2720), 
         .Z(n13568)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i3_4_lut_adj_551.init = 16'heca0;
    LUT4 i5183_4_lut (.A(n2713[10]), .B(n2775), .C(\address_7__N_549[1] ), 
         .D(spi_cmd[15]), .Z(n9976)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B)) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i5183_4_lut.init = 16'heece;
    LUT4 i28_4_lut (.A(n2713[11]), .B(n28723), .C(\address_7__N_549[1] ), 
         .D(n27596), .Z(n13_adj_6718)) /* synthesis lut_function=(A (B+((D)+!C))+!A (C (D))) */ ;   // c:/s_links/sources/spi_ctrl.v(16[45:52])
    defparam i28_4_lut.init = 16'hfa8a;
    LUT4 i22427_3_lut (.A(mem_rdata_update_N_729), .B(spi_cmd[15]), .C(spi_addr_valid_N_732), 
         .Z(n27596)) /* synthesis lut_function=(A+(B (C))) */ ;
    defparam i22427_3_lut.init = 16'heaea;
    LUT4 spi_cmd_start_reg_bdd_2_lut (.A(spi_csn_buf2_p), .B(spi_idle_N_747), 
         .Z(n28765)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam spi_cmd_start_reg_bdd_2_lut.init = 16'h2222;
    LUT4 i11_4_lut (.A(n2720), .B(wr_en), .C(mem_rdata_update_N_729), 
         .D(mem_wr), .Z(n7083)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i11_4_lut.init = 16'hcac0;
    LUT4 spi_cmd_start_reg_bdd_4_lut (.A(spi_cmd_start_reg_N_745), .B(spi_cmd_start_reg_N_746), 
         .C(spi_csn_buf2_p), .D(spi_idle_N_747), .Z(n28764)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+!(D))))) */ ;
    defparam spi_cmd_start_reg_bdd_4_lut.init = 16'h10f1;
    LUT4 mux_1736_i1_3_lut (.A(n13657), .B(\address_7__N_549[1] ), .C(spi_cmd_start_reg_N_746), 
         .Z(wr_en_N_697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam mux_1736_i1_3_lut.init = 16'hcaca;
    LUT4 i8762_4_lut (.A(n29186), .B(n29116), .C(n29241), .D(n7), .Z(n13657)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i8762_4_lut.init = 16'hc5c0;
    LUT4 i1_4_lut_adj_552 (.A(spi_cmd_start_reg_N_745), .B(n29240), .C(n8_adj_6709), 
         .D(n27630), .Z(n7)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i1_4_lut_adj_552.init = 16'hccdc;
    LUT4 mem_addr_2509_mux_6_i1_3_lut (.A(wb_dat_o[0]), .B(n37_adj_6725[0]), 
         .C(n7083), .Z(n47[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/spi_ctrl.v(382[42:54])
    defparam mem_addr_2509_mux_6_i1_3_lut.init = 16'hcaca;
    LUT4 i2182_2_lut (.A(spi_cmd_cnt), .B(n2724), .Z(spi_cmd_cnt_N_749)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/spi_ctrl.v(166[11] 390[18])
    defparam i2182_2_lut.init = 16'h6666;
    FD1P3AY spi_cmd_i0_i0_rep_593 (.D(wb_dat_o[0]), .SP(clk_enable_525), 
            .CK(clk), .Q(n29761)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=4, LSE_RCOL=21, LSE_LLINE=203, LSE_RLINE=225 */ ;   // c:/s_links/sources/spi_ctrl.v(159[17] 391[11])
    defparam spi_cmd_i0_i0_rep_593.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \quad_decoder(DEV_ID=5) 
//

module \quad_decoder(DEV_ID=5)  (quad_homing, n29220, pin_io_out_54, n95, 
            n66, n5647, n24, n32, quad_count, clk_1MHz, clk_1MHz_enable_171, 
            \spi_data_out_r_39__N_2104[0] , clk, \spi_data_out_r_39__N_2249[0] , 
            \quad_b[5] , quad_buffer, \mode[2]_derived_32 , clk_enable_28, 
            n29239, \spi_data_r[1] , n29762, clk_enable_131, \spi_data_r[0] , 
            \spi_data_r[31] , \spi_data_r[30] , \spi_data_r[29] , \spi_data_r[28] , 
            \spi_data_r[27] , \spi_data_r[26] , \spi_data_r[25] , \spi_data_r[24] , 
            \spi_data_r[23] , \spi_data_r[22] , \spi_data_r[21] , \spi_data_r[20] , 
            \spi_data_r[19] , \spi_data_r[18] , \spi_data_r[17] , \spi_data_r[16] , 
            \spi_data_r[15] , \spi_data_r[14] , \spi_data_r[13] , \spi_data_r[12] , 
            \spi_data_r[11] , \spi_data_r[10] , \spi_data_r[9] , \spi_data_r[8] , 
            \spi_data_r[7] , \spi_data_r[6] , \spi_data_r[5] , \spi_data_r[4] , 
            \spi_data_r[3] , \spi_data_r[2] , n29336, spi_data_out_r_39__N_2144, 
            spi_data_out_r_39__N_2332, quad_set_complete, quad_set_valid, 
            \quad_a[5] , \spi_data_out_r_39__N_2104[31] , \spi_data_out_r_39__N_2249[31] , 
            \spi_data_out_r_39__N_2104[30] , \spi_data_out_r_39__N_2249[30] , 
            \spi_data_out_r_39__N_2104[29] , \spi_data_out_r_39__N_2249[29] , 
            \spi_data_out_r_39__N_2104[28] , \spi_data_out_r_39__N_2249[28] , 
            \spi_data_out_r_39__N_2104[27] , \spi_data_out_r_39__N_2249[27] , 
            \spi_data_out_r_39__N_2104[26] , \spi_data_out_r_39__N_2249[26] , 
            \spi_data_out_r_39__N_2104[25] , \spi_data_out_r_39__N_2249[25] , 
            \spi_data_out_r_39__N_2104[24] , \spi_data_out_r_39__N_2249[24] , 
            \spi_data_out_r_39__N_2104[23] , \spi_data_out_r_39__N_2249[23] , 
            \spi_data_out_r_39__N_2104[22] , \spi_data_out_r_39__N_2249[22] , 
            \spi_data_out_r_39__N_2104[21] , \spi_data_out_r_39__N_2249[21] , 
            \spi_data_out_r_39__N_2104[20] , \spi_data_out_r_39__N_2249[20] , 
            \spi_data_out_r_39__N_2104[19] , \spi_data_out_r_39__N_2249[19] , 
            \spi_data_out_r_39__N_2104[18] , \spi_data_out_r_39__N_2249[18] , 
            \spi_data_out_r_39__N_2104[17] , \spi_data_out_r_39__N_2249[17] , 
            \spi_data_out_r_39__N_2104[16] , \spi_data_out_r_39__N_2249[16] , 
            \spi_data_out_r_39__N_2104[15] , \spi_data_out_r_39__N_2249[15] , 
            \spi_data_out_r_39__N_2104[14] , \spi_data_out_r_39__N_2249[14] , 
            \spi_data_out_r_39__N_2104[13] , \spi_data_out_r_39__N_2249[13] , 
            \spi_data_out_r_39__N_2104[12] , \spi_data_out_r_39__N_2249[12] , 
            \spi_data_out_r_39__N_2104[11] , \spi_data_out_r_39__N_2249[11] , 
            \spi_data_out_r_39__N_2104[10] , \spi_data_out_r_39__N_2249[10] , 
            \spi_data_out_r_39__N_2104[9] , \spi_data_out_r_39__N_2249[9] , 
            \spi_data_out_r_39__N_2104[8] , \spi_data_out_r_39__N_2249[8] , 
            \spi_data_out_r_39__N_2104[7] , \spi_data_out_r_39__N_2249[7] , 
            \spi_data_out_r_39__N_2104[6] , \spi_data_out_r_39__N_2249[6] , 
            \spi_data_out_r_39__N_2104[5] , \spi_data_out_r_39__N_2249[5] , 
            \spi_data_out_r_39__N_2104[4] , \spi_data_out_r_39__N_2249[4] , 
            \spi_data_out_r_39__N_2104[3] , \spi_data_out_r_39__N_2249[3] , 
            \spi_data_out_r_39__N_2104[2] , \spi_data_out_r_39__N_2249[2] , 
            \spi_data_out_r_39__N_2104[1] , \spi_data_out_r_39__N_2249[1] , 
            resetn_c, GND_net, clk_enable_519, n29079, n21446) /* synthesis syn_module_defined=1 */ ;
    output [1:0]quad_homing;
    input n29220;
    input pin_io_out_54;
    output n95;
    output n66;
    input n5647;
    input n24;
    output n32;
    output [31:0]quad_count;
    input clk_1MHz;
    input clk_1MHz_enable_171;
    output \spi_data_out_r_39__N_2104[0] ;
    input clk;
    input \spi_data_out_r_39__N_2249[0] ;
    input \quad_b[5] ;
    output [31:0]quad_buffer;
    input \mode[2]_derived_32 ;
    input clk_enable_28;
    input n29239;
    input \spi_data_r[1] ;
    input n29762;
    input clk_enable_131;
    input \spi_data_r[0] ;
    input \spi_data_r[31] ;
    input \spi_data_r[30] ;
    input \spi_data_r[29] ;
    input \spi_data_r[28] ;
    input \spi_data_r[27] ;
    input \spi_data_r[26] ;
    input \spi_data_r[25] ;
    input \spi_data_r[24] ;
    input \spi_data_r[23] ;
    input \spi_data_r[22] ;
    input \spi_data_r[21] ;
    input \spi_data_r[20] ;
    input \spi_data_r[19] ;
    input \spi_data_r[18] ;
    input \spi_data_r[17] ;
    input \spi_data_r[16] ;
    input \spi_data_r[15] ;
    input \spi_data_r[14] ;
    input \spi_data_r[13] ;
    input \spi_data_r[12] ;
    input \spi_data_r[11] ;
    input \spi_data_r[10] ;
    input \spi_data_r[9] ;
    input \spi_data_r[8] ;
    input \spi_data_r[7] ;
    input \spi_data_r[6] ;
    input \spi_data_r[5] ;
    input \spi_data_r[4] ;
    input \spi_data_r[3] ;
    input \spi_data_r[2] ;
    output n29336;
    output spi_data_out_r_39__N_2144;
    input spi_data_out_r_39__N_2332;
    output quad_set_complete;
    output quad_set_valid;
    input \quad_a[5] ;
    output \spi_data_out_r_39__N_2104[31] ;
    input \spi_data_out_r_39__N_2249[31] ;
    output \spi_data_out_r_39__N_2104[30] ;
    input \spi_data_out_r_39__N_2249[30] ;
    output \spi_data_out_r_39__N_2104[29] ;
    input \spi_data_out_r_39__N_2249[29] ;
    output \spi_data_out_r_39__N_2104[28] ;
    input \spi_data_out_r_39__N_2249[28] ;
    output \spi_data_out_r_39__N_2104[27] ;
    input \spi_data_out_r_39__N_2249[27] ;
    output \spi_data_out_r_39__N_2104[26] ;
    input \spi_data_out_r_39__N_2249[26] ;
    output \spi_data_out_r_39__N_2104[25] ;
    input \spi_data_out_r_39__N_2249[25] ;
    output \spi_data_out_r_39__N_2104[24] ;
    input \spi_data_out_r_39__N_2249[24] ;
    output \spi_data_out_r_39__N_2104[23] ;
    input \spi_data_out_r_39__N_2249[23] ;
    output \spi_data_out_r_39__N_2104[22] ;
    input \spi_data_out_r_39__N_2249[22] ;
    output \spi_data_out_r_39__N_2104[21] ;
    input \spi_data_out_r_39__N_2249[21] ;
    output \spi_data_out_r_39__N_2104[20] ;
    input \spi_data_out_r_39__N_2249[20] ;
    output \spi_data_out_r_39__N_2104[19] ;
    input \spi_data_out_r_39__N_2249[19] ;
    output \spi_data_out_r_39__N_2104[18] ;
    input \spi_data_out_r_39__N_2249[18] ;
    output \spi_data_out_r_39__N_2104[17] ;
    input \spi_data_out_r_39__N_2249[17] ;
    output \spi_data_out_r_39__N_2104[16] ;
    input \spi_data_out_r_39__N_2249[16] ;
    output \spi_data_out_r_39__N_2104[15] ;
    input \spi_data_out_r_39__N_2249[15] ;
    output \spi_data_out_r_39__N_2104[14] ;
    input \spi_data_out_r_39__N_2249[14] ;
    output \spi_data_out_r_39__N_2104[13] ;
    input \spi_data_out_r_39__N_2249[13] ;
    output \spi_data_out_r_39__N_2104[12] ;
    input \spi_data_out_r_39__N_2249[12] ;
    output \spi_data_out_r_39__N_2104[11] ;
    input \spi_data_out_r_39__N_2249[11] ;
    output \spi_data_out_r_39__N_2104[10] ;
    input \spi_data_out_r_39__N_2249[10] ;
    output \spi_data_out_r_39__N_2104[9] ;
    input \spi_data_out_r_39__N_2249[9] ;
    output \spi_data_out_r_39__N_2104[8] ;
    input \spi_data_out_r_39__N_2249[8] ;
    output \spi_data_out_r_39__N_2104[7] ;
    input \spi_data_out_r_39__N_2249[7] ;
    output \spi_data_out_r_39__N_2104[6] ;
    input \spi_data_out_r_39__N_2249[6] ;
    output \spi_data_out_r_39__N_2104[5] ;
    input \spi_data_out_r_39__N_2249[5] ;
    output \spi_data_out_r_39__N_2104[4] ;
    input \spi_data_out_r_39__N_2249[4] ;
    output \spi_data_out_r_39__N_2104[3] ;
    input \spi_data_out_r_39__N_2249[3] ;
    output \spi_data_out_r_39__N_2104[2] ;
    input \spi_data_out_r_39__N_2249[2] ;
    output \spi_data_out_r_39__N_2104[1] ;
    input \spi_data_out_r_39__N_2249[1] ;
    input resetn_c;
    input GND_net;
    input clk_enable_519;
    input n29079;
    output n21446;
    
    wire [1:0]AB /* synthesis ASYNC_REG="TRUE" */ ;   // c:/s_links/sources/quad_decoder.v(106[36:38])
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire [1:0]sync /* synthesis ASYNC_REG="TRUE" */ ;   // c:/s_links/sources/quad_decoder.v(106[30:34])
    wire \mode[2]_derived_32  /* synthesis is_clock=1, SET_AS_NETWORK=\stepper_ins[5].u_stepper/mode[2]_derived_32 */ ;   // c:/s_links/sources/slot_cards/stepper.v(53[11:15])
    wire [31:0]n6171;
    wire [31:0]quad_set;   // c:/s_links/sources/quad_decoder.v(40[31:39])
    
    wire n10788, n10786, n29221, n10784, n10782, n29222;
    wire [3:0]n2281;
    
    wire n4, n9596, n6, n26889, n9956, n10780, n10778, n10776, 
        n10774, n10772, n10770, n10768, n10766, n10764, n29004, 
        n10762, n29323, n29324, n29325, n10760, n21498, n21501, 
        n10758, n10756, n10754, n10752, n10750, n10748, n10746, 
        n10744, n10742, n10740, n10738, n10736, n10734, n10732, 
        n10792, n10790, n25130, n25129, n25128, n25127, n25126, 
        n25125, n25124, n25123, n25122, n25121, n25120, n25119, 
        n25118, n25117, n25116, n25115;
    
    LUT4 i109_2_lut_3_lut_4_lut (.A(quad_homing[0]), .B(quad_homing[1]), 
         .C(n29220), .D(pin_io_out_54), .Z(n95)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam i109_2_lut_3_lut_4_lut.init = 16'hfdff;
    LUT4 i1_2_lut_3_lut_4_lut (.A(quad_homing[0]), .B(quad_homing[1]), .C(n29220), 
         .D(pin_io_out_54), .Z(n66)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0200;
    LUT4 i5995_4_lut (.A(n6171[29]), .B(quad_set[29]), .C(n5647), .D(n24), 
         .Z(n10788)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5995_4_lut.init = 16'hc0ca;
    LUT4 i5993_4_lut (.A(n6171[28]), .B(quad_set[28]), .C(n5647), .D(n24), 
         .Z(n10786)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5993_4_lut.init = 16'hc0ca;
    LUT4 i35_2_lut_rep_493 (.A(AB[1]), .B(AB[0]), .Z(n29221)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/s_links/sources/quad_decoder.v(106[36:38])
    defparam i35_2_lut_rep_493.init = 16'h6666;
    LUT4 i5991_4_lut (.A(n6171[27]), .B(quad_set[27]), .C(n5647), .D(n24), 
         .Z(n10784)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5991_4_lut.init = 16'hc0ca;
    LUT4 i5989_4_lut (.A(n6171[26]), .B(quad_set[26]), .C(n5647), .D(n24), 
         .Z(n10782)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5989_4_lut.init = 16'hc0ca;
    LUT4 i46_4_lut_3_lut_4_lut (.A(AB[1]), .B(AB[0]), .C(n29222), .D(n2281[3]), 
         .Z(n32)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B !((D)+!C))) */ ;   // c:/s_links/sources/quad_decoder.v(106[36:38])
    defparam i46_4_lut_3_lut_4_lut.init = 16'h9969;
    LUT4 i16576_4_lut_4_lut (.A(AB[1]), .B(AB[0]), .C(n4), .D(n2281[3]), 
         .Z(n9596)) /* synthesis lut_function=(A (B (C+(D)))+!A !(B ((D)+!C)+!B !(D))) */ ;   // c:/s_links/sources/quad_decoder.v(106[36:38])
    defparam i16576_4_lut_4_lut.init = 16'h99c0;
    LUT4 i1_4_lut_4_lut (.A(AB[1]), .B(AB[0]), .C(n2281[1]), .D(n6), 
         .Z(n26889)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C+(D))))) */ ;   // c:/s_links/sources/quad_decoder.v(106[36:38])
    defparam i1_4_lut_4_lut.init = 16'h6460;
    LUT4 i22403_2_lut_rep_494 (.A(n2281[1]), .B(n2281[2]), .Z(n29222)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i22403_2_lut_rep_494.init = 16'heeee;
    FD1P3AX quad_count_i0_i0 (.D(n9956), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i0.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut (.A(n2281[1]), .B(n2281[2]), .C(AB[1]), .Z(n4)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'he0e0;
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_2249[0] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX sync_i0 (.D(\quad_b[5] ), .CK(clk_1MHz), .Q(sync[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam sync_i0.GSR = "DISABLED";
    LUT4 i5987_4_lut (.A(n6171[25]), .B(quad_set[25]), .C(n5647), .D(n24), 
         .Z(n10780)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5987_4_lut.init = 16'hc0ca;
    FD1S3AX AB_i0 (.D(sync[0]), .CK(clk_1MHz), .Q(AB[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam AB_i0.GSR = "DISABLED";
    FD1S3AX quad_buffer_i0 (.D(quad_count[0]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i0.GSR = "DISABLED";
    LUT4 i5985_4_lut (.A(n6171[24]), .B(quad_set[24]), .C(n5647), .D(n24), 
         .Z(n10778)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5985_4_lut.init = 16'hc0ca;
    LUT4 i5983_4_lut (.A(n6171[23]), .B(quad_set[23]), .C(n5647), .D(n24), 
         .Z(n10776)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5983_4_lut.init = 16'hc0ca;
    FD1P3IX quad_homing__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_28), .CD(n29239), 
            .CK(clk), .Q(quad_homing[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam quad_homing__i1.GSR = "DISABLED";
    LUT4 i5981_4_lut (.A(n6171[22]), .B(quad_set[22]), .C(n5647), .D(n24), 
         .Z(n10774)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5981_4_lut.init = 16'hc0ca;
    LUT4 i5979_4_lut (.A(n6171[21]), .B(quad_set[21]), .C(n5647), .D(n24), 
         .Z(n10772)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5979_4_lut.init = 16'hc0ca;
    LUT4 i5977_4_lut (.A(n6171[20]), .B(quad_set[20]), .C(n5647), .D(n24), 
         .Z(n10770)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5977_4_lut.init = 16'hc0ca;
    LUT4 i5975_4_lut (.A(n6171[19]), .B(quad_set[19]), .C(n5647), .D(n24), 
         .Z(n10768)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5975_4_lut.init = 16'hc0ca;
    LUT4 i5973_4_lut (.A(n6171[18]), .B(quad_set[18]), .C(n5647), .D(n24), 
         .Z(n10766)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5973_4_lut.init = 16'hc0ca;
    FD1P3IX quad_homing__i0 (.D(n29762), .SP(clk_enable_28), .CD(n29239), 
            .CK(clk), .Q(quad_homing[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(65[8] 72[4])
    defparam quad_homing__i0.GSR = "DISABLED";
    FD1P3IX quad_set__i0 (.D(\spi_data_r[0] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i0.GSR = "DISABLED";
    LUT4 i5971_4_lut (.A(n6171[17]), .B(quad_set[17]), .C(n5647), .D(n24), 
         .Z(n10764)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5971_4_lut.init = 16'hc0ca;
    FD1S3JX state_FSM_i0 (.D(n29004), .CK(clk_1MHz), .PD(n29239), .Q(n2281[0]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i0.GSR = "DISABLED";
    LUT4 i5969_4_lut (.A(n6171[16]), .B(quad_set[16]), .C(n5647), .D(n24), 
         .Z(n10762)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5969_4_lut.init = 16'hc0ca;
    PFUMX i23158 (.BLUT(n29323), .ALUT(n29324), .C0(n2281[3]), .Z(n29325));
    FD1P3IX quad_set__i31 (.D(\spi_data_r[31] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i31.GSR = "DISABLED";
    FD1P3IX quad_set__i30 (.D(\spi_data_r[30] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i30.GSR = "DISABLED";
    FD1P3IX quad_set__i29 (.D(\spi_data_r[29] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i29.GSR = "DISABLED";
    FD1P3IX quad_set__i28 (.D(\spi_data_r[28] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i28.GSR = "DISABLED";
    FD1P3IX quad_set__i27 (.D(\spi_data_r[27] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i27.GSR = "DISABLED";
    FD1P3IX quad_set__i26 (.D(\spi_data_r[26] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i26.GSR = "DISABLED";
    FD1P3IX quad_set__i25 (.D(\spi_data_r[25] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i25.GSR = "DISABLED";
    FD1P3IX quad_set__i24 (.D(\spi_data_r[24] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i24.GSR = "DISABLED";
    FD1P3IX quad_set__i23 (.D(\spi_data_r[23] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i23.GSR = "DISABLED";
    FD1P3IX quad_set__i22 (.D(\spi_data_r[22] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i22.GSR = "DISABLED";
    FD1P3IX quad_set__i21 (.D(\spi_data_r[21] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i21.GSR = "DISABLED";
    FD1P3IX quad_set__i20 (.D(\spi_data_r[20] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i20.GSR = "DISABLED";
    FD1P3IX quad_set__i19 (.D(\spi_data_r[19] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i19.GSR = "DISABLED";
    FD1P3IX quad_set__i18 (.D(\spi_data_r[18] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i18.GSR = "DISABLED";
    FD1P3IX quad_set__i17 (.D(\spi_data_r[17] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i17.GSR = "DISABLED";
    FD1P3IX quad_set__i16 (.D(\spi_data_r[16] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i16.GSR = "DISABLED";
    FD1P3IX quad_set__i15 (.D(\spi_data_r[15] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i15.GSR = "DISABLED";
    FD1P3IX quad_set__i14 (.D(\spi_data_r[14] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i14.GSR = "DISABLED";
    FD1P3IX quad_set__i13 (.D(\spi_data_r[13] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i13.GSR = "DISABLED";
    FD1P3IX quad_set__i12 (.D(\spi_data_r[12] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i12.GSR = "DISABLED";
    FD1P3IX quad_set__i11 (.D(\spi_data_r[11] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i11.GSR = "DISABLED";
    FD1P3IX quad_set__i10 (.D(\spi_data_r[10] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i10.GSR = "DISABLED";
    FD1P3IX quad_set__i9 (.D(\spi_data_r[9] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i9.GSR = "DISABLED";
    FD1P3IX quad_set__i8 (.D(\spi_data_r[8] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i8.GSR = "DISABLED";
    FD1P3IX quad_set__i7 (.D(\spi_data_r[7] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i7.GSR = "DISABLED";
    FD1P3IX quad_set__i6 (.D(\spi_data_r[6] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i6.GSR = "DISABLED";
    FD1P3IX quad_set__i5 (.D(\spi_data_r[5] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i5.GSR = "DISABLED";
    FD1P3IX quad_set__i4 (.D(\spi_data_r[4] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i4.GSR = "DISABLED";
    FD1P3IX quad_set__i3 (.D(\spi_data_r[3] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i3.GSR = "DISABLED";
    FD1P3IX quad_set__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i2.GSR = "DISABLED";
    FD1P3IX quad_set__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_131), .CD(n29239), 
            .CK(clk), .Q(quad_set[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set__i1.GSR = "DISABLED";
    LUT4 i5967_4_lut (.A(n6171[15]), .B(quad_set[15]), .C(n5647), .D(n24), 
         .Z(n10760)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5967_4_lut.init = 16'hc0ca;
    LUT4 i16563_3_lut_4_lut (.A(AB[1]), .B(AB[0]), .C(n2281[3]), .D(n21498), 
         .Z(n21501)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam i16563_3_lut_4_lut.init = 16'h2f20;
    LUT4 i5965_4_lut (.A(n6171[14]), .B(quad_set[14]), .C(n5647), .D(n24), 
         .Z(n10758)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5965_4_lut.init = 16'hc0ca;
    LUT4 i5963_4_lut (.A(n6171[13]), .B(quad_set[13]), .C(n5647), .D(n24), 
         .Z(n10756)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5963_4_lut.init = 16'hc0ca;
    LUT4 n2282_bdd_4_lut_23171 (.A(n2281[3]), .B(n29222), .C(AB[0]), .D(AB[1]), 
         .Z(n29336)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam n2282_bdd_4_lut_23171.init = 16'hb44b;
    LUT4 i5961_4_lut (.A(n6171[12]), .B(quad_set[12]), .C(n5647), .D(n24), 
         .Z(n10754)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5961_4_lut.init = 16'hc0ca;
    FD1S3IX i41_407 (.D(spi_data_out_r_39__N_2332), .CK(clk), .CD(n29239), 
            .Q(spi_data_out_r_39__N_2144)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam i41_407.GSR = "DISABLED";
    LUT4 i5959_4_lut (.A(n6171[11]), .B(quad_set[11]), .C(n5647), .D(n24), 
         .Z(n10752)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5959_4_lut.init = 16'hc0ca;
    FD1S3IX quad_set_complete_451 (.D(quad_set_valid), .CK(clk_1MHz), .CD(n29239), 
            .Q(quad_set_complete)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_set_complete_451.GSR = "DISABLED";
    LUT4 i5957_4_lut (.A(n6171[10]), .B(quad_set[10]), .C(n5647), .D(n24), 
         .Z(n10750)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5957_4_lut.init = 16'hc0ca;
    LUT4 i5955_4_lut (.A(n6171[9]), .B(quad_set[9]), .C(n5647), .D(n24), 
         .Z(n10748)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5955_4_lut.init = 16'hc0ca;
    LUT4 i5953_4_lut (.A(n6171[8]), .B(quad_set[8]), .C(n5647), .D(n24), 
         .Z(n10746)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5953_4_lut.init = 16'hc0ca;
    LUT4 i5951_4_lut (.A(n6171[7]), .B(quad_set[7]), .C(n5647), .D(n24), 
         .Z(n10744)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5951_4_lut.init = 16'hc0ca;
    LUT4 i5949_4_lut (.A(n6171[6]), .B(quad_set[6]), .C(n5647), .D(n24), 
         .Z(n10742)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5949_4_lut.init = 16'hc0ca;
    LUT4 i5947_4_lut (.A(n6171[5]), .B(quad_set[5]), .C(n5647), .D(n24), 
         .Z(n10740)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5947_4_lut.init = 16'hc0ca;
    LUT4 n2285_bdd_4_lut (.A(n2281[0]), .B(n29222), .C(AB[1]), .D(AB[0]), 
         .Z(n29004)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !((C+(D))+!B)) */ ;
    defparam n2285_bdd_4_lut.init = 16'ha00e;
    LUT4 i5945_4_lut (.A(n6171[4]), .B(quad_set[4]), .C(n5647), .D(n24), 
         .Z(n10738)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5945_4_lut.init = 16'hc0ca;
    LUT4 i5943_4_lut (.A(n6171[3]), .B(quad_set[3]), .C(n5647), .D(n24), 
         .Z(n10736)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5943_4_lut.init = 16'hc0ca;
    LUT4 i5941_4_lut (.A(n6171[2]), .B(quad_set[2]), .C(n5647), .D(n24), 
         .Z(n10734)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5941_4_lut.init = 16'hc0ca;
    LUT4 i5939_4_lut (.A(n6171[1]), .B(quad_set[1]), .C(n5647), .D(n24), 
         .Z(n10732)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5939_4_lut.init = 16'hc0ca;
    FD1S3AX quad_buffer_i31 (.D(quad_count[31]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i31.GSR = "DISABLED";
    FD1S3AX quad_buffer_i30 (.D(quad_count[30]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i30.GSR = "DISABLED";
    FD1S3AX quad_buffer_i29 (.D(quad_count[29]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i29.GSR = "DISABLED";
    FD1S3AX quad_buffer_i28 (.D(quad_count[28]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i28.GSR = "DISABLED";
    FD1S3AX quad_buffer_i27 (.D(quad_count[27]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i27.GSR = "DISABLED";
    FD1S3AX quad_buffer_i26 (.D(quad_count[26]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i26.GSR = "DISABLED";
    FD1S3AX quad_buffer_i25 (.D(quad_count[25]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i25.GSR = "DISABLED";
    FD1S3AX quad_buffer_i24 (.D(quad_count[24]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i24.GSR = "DISABLED";
    FD1S3AX quad_buffer_i23 (.D(quad_count[23]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i23.GSR = "DISABLED";
    FD1S3AX quad_buffer_i22 (.D(quad_count[22]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i22.GSR = "DISABLED";
    FD1S3AX quad_buffer_i21 (.D(quad_count[21]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i21.GSR = "DISABLED";
    FD1S3AX quad_buffer_i20 (.D(quad_count[20]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i20.GSR = "DISABLED";
    FD1S3AX quad_buffer_i19 (.D(quad_count[19]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i19.GSR = "DISABLED";
    FD1S3AX quad_buffer_i18 (.D(quad_count[18]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i18.GSR = "DISABLED";
    FD1S3AX quad_buffer_i17 (.D(quad_count[17]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i17.GSR = "DISABLED";
    FD1S3AX quad_buffer_i16 (.D(quad_count[16]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i16.GSR = "DISABLED";
    FD1S3AX quad_buffer_i15 (.D(quad_count[15]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i15.GSR = "DISABLED";
    FD1S3AX quad_buffer_i14 (.D(quad_count[14]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i14.GSR = "DISABLED";
    FD1S3AX quad_buffer_i13 (.D(quad_count[13]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i13.GSR = "DISABLED";
    FD1S3AX quad_buffer_i12 (.D(quad_count[12]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i12.GSR = "DISABLED";
    FD1S3AX quad_buffer_i11 (.D(quad_count[11]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i11.GSR = "DISABLED";
    FD1S3AX quad_buffer_i10 (.D(quad_count[10]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i10.GSR = "DISABLED";
    FD1S3AX quad_buffer_i9 (.D(quad_count[9]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i9.GSR = "DISABLED";
    FD1S3AX quad_buffer_i8 (.D(quad_count[8]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i8.GSR = "DISABLED";
    FD1S3AX quad_buffer_i7 (.D(quad_count[7]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i7.GSR = "DISABLED";
    FD1S3AX quad_buffer_i6 (.D(quad_count[6]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i6.GSR = "DISABLED";
    FD1S3AX quad_buffer_i5 (.D(quad_count[5]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i5.GSR = "DISABLED";
    FD1S3AX quad_buffer_i4 (.D(quad_count[4]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i4.GSR = "DISABLED";
    FD1S3AX quad_buffer_i3 (.D(quad_count[3]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i3.GSR = "DISABLED";
    FD1S3AX quad_buffer_i2 (.D(quad_count[2]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i2.GSR = "DISABLED";
    FD1S3AX quad_buffer_i1 (.D(quad_count[1]), .CK(\mode[2]_derived_32 ), 
            .Q(quad_buffer[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(214[8] 216[4])
    defparam quad_buffer_i1.GSR = "DISABLED";
    FD1S3AX AB_i1 (.D(sync[1]), .CK(clk_1MHz), .Q(AB[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam AB_i1.GSR = "DISABLED";
    FD1S3AX sync_i1 (.D(\quad_a[5] ), .CK(clk_1MHz), .Q(sync[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(110[8] 114[4])
    defparam sync_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_2249[31] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[31] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i31 (.D(\spi_data_out_r_39__N_2249[30] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[30] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i30 (.D(\spi_data_out_r_39__N_2249[29] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i29 (.D(\spi_data_out_r_39__N_2249[28] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i28 (.D(\spi_data_out_r_39__N_2249[27] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i27 (.D(\spi_data_out_r_39__N_2249[26] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i26 (.D(\spi_data_out_r_39__N_2249[25] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i25 (.D(\spi_data_out_r_39__N_2249[24] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i24 (.D(\spi_data_out_r_39__N_2249[23] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i23 (.D(\spi_data_out_r_39__N_2249[22] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i22 (.D(\spi_data_out_r_39__N_2249[21] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i21 (.D(\spi_data_out_r_39__N_2249[20] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i20 (.D(\spi_data_out_r_39__N_2249[19] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i19 (.D(\spi_data_out_r_39__N_2249[18] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i18 (.D(\spi_data_out_r_39__N_2249[17] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i17 (.D(\spi_data_out_r_39__N_2249[16] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i16 (.D(\spi_data_out_r_39__N_2249[15] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_2249[14] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_2249[13] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_2249[12] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_2249[11] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_2249[10] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_2249[9] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_2249[8] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_2249[7] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_2249[6] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_2249[5] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_2249[4] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_2249[3] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_2249[2] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_2249[1] ), .CK(clk), 
            .Q(\spi_data_out_r_39__N_2104[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(75[8] 84[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    LUT4 i16560_4_lut (.A(AB[0]), .B(AB[1]), .C(n2281[2]), .D(n2281[1]), 
         .Z(n21498)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C+(D)))+!A (B+!(C)))) */ ;
    defparam i16560_4_lut.init = 16'h1812;
    FD1P3AX quad_count_i0_i31 (.D(n10792), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i31.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i30 (.D(n10790), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i30.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i29 (.D(n10788), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i29.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i28 (.D(n10786), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i28.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i27 (.D(n10784), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i27.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i26 (.D(n10782), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i26.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i25 (.D(n10780), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i25.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i24 (.D(n10778), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i24.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i23 (.D(n10776), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i23.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i22 (.D(n10774), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i22.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i21 (.D(n10772), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i21.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i20 (.D(n10770), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i20.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i19 (.D(n10768), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i19.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i18 (.D(n10766), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i18.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i17 (.D(n10764), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i17.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i16 (.D(n10762), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i16.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i15 (.D(n10760), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i15.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i14 (.D(n10758), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i14.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i13 (.D(n10756), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i13.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i12 (.D(n10754), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i12.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i11 (.D(n10752), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i11.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i10 (.D(n10750), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i10.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i9 (.D(n10748), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i9.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i8 (.D(n10746), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i8.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i7 (.D(n10744), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i7.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i6 (.D(n10742), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i6.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i5 (.D(n10740), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i5.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i4 (.D(n10738), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i4.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i3 (.D(n10736), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i3.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i2 (.D(n10734), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i2.GSR = "DISABLED";
    FD1P3AX quad_count_i0_i1 (.D(n10732), .SP(clk_1MHz_enable_171), .CK(clk_1MHz), 
            .Q(quad_count[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(118[8] 169[4])
    defparam quad_count_i0_i1.GSR = "DISABLED";
    LUT4 i5999_4_lut (.A(n6171[31]), .B(quad_set[31]), .C(n5647), .D(n24), 
         .Z(n10792)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5999_4_lut.init = 16'hc0ca;
    LUT4 i5997_4_lut (.A(n6171[30]), .B(quad_set[30]), .C(n5647), .D(n24), 
         .Z(n10790)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5997_4_lut.init = 16'hc0ca;
    LUT4 i33_4_lut_then_3_lut (.A(n2281[2]), .B(AB[0]), .C(AB[1]), .Z(n29324)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;
    defparam i33_4_lut_then_3_lut.init = 16'h3838;
    FD1S3IX state_FSM_i1 (.D(n26889), .CK(clk_1MHz), .CD(n29239), .Q(n2281[1]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i1.GSR = "DISABLED";
    FD1S3IX state_FSM_i2 (.D(n29325), .CK(clk_1MHz), .CD(n29239), .Q(n2281[2]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i2.GSR = "DISABLED";
    FD1S3IX state_FSM_i3 (.D(n9596), .CK(clk_1MHz), .CD(n29239), .Q(n2281[3]));   // c:/s_links/sources/quad_decoder.v(137[4] 166[12])
    defparam state_FSM_i3.GSR = "DISABLED";
    CCU2D add_1980_33 (.A0(resetn_c), .B0(n21501), .C0(quad_count[30]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[31]), 
          .D1(GND_net), .CIN(n25130), .S0(n6171[30]), .S1(n6171[31]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_33.INIT0 = 16'h7878;
    defparam add_1980_33.INIT1 = 16'h7878;
    defparam add_1980_33.INJECT1_0 = "NO";
    defparam add_1980_33.INJECT1_1 = "NO";
    CCU2D add_1980_31 (.A0(resetn_c), .B0(n21501), .C0(quad_count[28]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[29]), 
          .D1(GND_net), .CIN(n25129), .COUT(n25130), .S0(n6171[28]), 
          .S1(n6171[29]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_31.INIT0 = 16'h7878;
    defparam add_1980_31.INIT1 = 16'h7878;
    defparam add_1980_31.INJECT1_0 = "NO";
    defparam add_1980_31.INJECT1_1 = "NO";
    CCU2D add_1980_29 (.A0(resetn_c), .B0(n21501), .C0(quad_count[26]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[27]), 
          .D1(GND_net), .CIN(n25128), .COUT(n25129), .S0(n6171[26]), 
          .S1(n6171[27]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_29.INIT0 = 16'h7878;
    defparam add_1980_29.INIT1 = 16'h7878;
    defparam add_1980_29.INJECT1_0 = "NO";
    defparam add_1980_29.INJECT1_1 = "NO";
    CCU2D add_1980_27 (.A0(resetn_c), .B0(n21501), .C0(quad_count[24]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[25]), 
          .D1(GND_net), .CIN(n25127), .COUT(n25128), .S0(n6171[24]), 
          .S1(n6171[25]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_27.INIT0 = 16'h7878;
    defparam add_1980_27.INIT1 = 16'h7878;
    defparam add_1980_27.INJECT1_0 = "NO";
    defparam add_1980_27.INJECT1_1 = "NO";
    CCU2D add_1980_25 (.A0(resetn_c), .B0(n21501), .C0(quad_count[22]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[23]), 
          .D1(GND_net), .CIN(n25126), .COUT(n25127), .S0(n6171[22]), 
          .S1(n6171[23]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_25.INIT0 = 16'h7878;
    defparam add_1980_25.INIT1 = 16'h7878;
    defparam add_1980_25.INJECT1_0 = "NO";
    defparam add_1980_25.INJECT1_1 = "NO";
    CCU2D add_1980_23 (.A0(resetn_c), .B0(n21501), .C0(quad_count[20]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[21]), 
          .D1(GND_net), .CIN(n25125), .COUT(n25126), .S0(n6171[20]), 
          .S1(n6171[21]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_23.INIT0 = 16'h7878;
    defparam add_1980_23.INIT1 = 16'h7878;
    defparam add_1980_23.INJECT1_0 = "NO";
    defparam add_1980_23.INJECT1_1 = "NO";
    CCU2D add_1980_21 (.A0(resetn_c), .B0(n21501), .C0(quad_count[18]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[19]), 
          .D1(GND_net), .CIN(n25124), .COUT(n25125), .S0(n6171[18]), 
          .S1(n6171[19]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_21.INIT0 = 16'h7878;
    defparam add_1980_21.INIT1 = 16'h7878;
    defparam add_1980_21.INJECT1_0 = "NO";
    defparam add_1980_21.INJECT1_1 = "NO";
    CCU2D add_1980_19 (.A0(resetn_c), .B0(n21501), .C0(quad_count[16]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[17]), 
          .D1(GND_net), .CIN(n25123), .COUT(n25124), .S0(n6171[16]), 
          .S1(n6171[17]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_19.INIT0 = 16'h7878;
    defparam add_1980_19.INIT1 = 16'h7878;
    defparam add_1980_19.INJECT1_0 = "NO";
    defparam add_1980_19.INJECT1_1 = "NO";
    CCU2D add_1980_17 (.A0(resetn_c), .B0(n21501), .C0(quad_count[14]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[15]), 
          .D1(GND_net), .CIN(n25122), .COUT(n25123), .S0(n6171[14]), 
          .S1(n6171[15]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_17.INIT0 = 16'h7878;
    defparam add_1980_17.INIT1 = 16'h7878;
    defparam add_1980_17.INJECT1_0 = "NO";
    defparam add_1980_17.INJECT1_1 = "NO";
    LUT4 i1_3_lut (.A(n2281[3]), .B(n2281[1]), .C(n2281[0]), .Z(n6)) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam i1_3_lut.init = 16'hbaba;
    CCU2D add_1980_15 (.A0(resetn_c), .B0(n21501), .C0(quad_count[12]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[13]), 
          .D1(GND_net), .CIN(n25121), .COUT(n25122), .S0(n6171[12]), 
          .S1(n6171[13]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_15.INIT0 = 16'h7878;
    defparam add_1980_15.INIT1 = 16'h7878;
    defparam add_1980_15.INJECT1_0 = "NO";
    defparam add_1980_15.INJECT1_1 = "NO";
    CCU2D add_1980_13 (.A0(resetn_c), .B0(n21501), .C0(quad_count[10]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[11]), 
          .D1(GND_net), .CIN(n25120), .COUT(n25121), .S0(n6171[10]), 
          .S1(n6171[11]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_13.INIT0 = 16'h7878;
    defparam add_1980_13.INIT1 = 16'h7878;
    defparam add_1980_13.INJECT1_0 = "NO";
    defparam add_1980_13.INJECT1_1 = "NO";
    CCU2D add_1980_11 (.A0(resetn_c), .B0(n21501), .C0(quad_count[8]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[9]), 
          .D1(GND_net), .CIN(n25119), .COUT(n25120), .S0(n6171[8]), 
          .S1(n6171[9]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_11.INIT0 = 16'h7878;
    defparam add_1980_11.INIT1 = 16'h7878;
    defparam add_1980_11.INJECT1_0 = "NO";
    defparam add_1980_11.INJECT1_1 = "NO";
    CCU2D add_1980_9 (.A0(resetn_c), .B0(n21501), .C0(quad_count[6]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[7]), 
          .D1(GND_net), .CIN(n25118), .COUT(n25119), .S0(n6171[6]), 
          .S1(n6171[7]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_9.INIT0 = 16'h7878;
    defparam add_1980_9.INIT1 = 16'h7878;
    defparam add_1980_9.INJECT1_0 = "NO";
    defparam add_1980_9.INJECT1_1 = "NO";
    CCU2D add_1980_7 (.A0(resetn_c), .B0(n21501), .C0(quad_count[4]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[5]), 
          .D1(GND_net), .CIN(n25117), .COUT(n25118), .S0(n6171[4]), 
          .S1(n6171[5]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_7.INIT0 = 16'h7878;
    defparam add_1980_7.INIT1 = 16'h7878;
    defparam add_1980_7.INJECT1_0 = "NO";
    defparam add_1980_7.INJECT1_1 = "NO";
    CCU2D add_1980_5 (.A0(resetn_c), .B0(n21501), .C0(quad_count[2]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[3]), 
          .D1(GND_net), .CIN(n25116), .COUT(n25117), .S0(n6171[2]), 
          .S1(n6171[3]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_5.INIT0 = 16'h7878;
    defparam add_1980_5.INIT1 = 16'h7878;
    defparam add_1980_5.INJECT1_0 = "NO";
    defparam add_1980_5.INJECT1_1 = "NO";
    LUT4 i33_4_lut_else_3_lut (.A(n2281[2]), .B(AB[0]), .C(AB[1]), .D(n2281[0]), 
         .Z(n29323)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C (D))))) */ ;
    defparam i33_4_lut_else_3_lut.init = 16'h3828;
    CCU2D add_1980_3 (.A0(resetn_c), .B0(n21501), .C0(quad_count[0]), 
          .D0(GND_net), .A1(resetn_c), .B1(n21501), .C1(quad_count[1]), 
          .D1(GND_net), .CIN(n25115), .COUT(n25116), .S0(n6171[0]), 
          .S1(n6171[1]));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_3.INIT0 = 16'h8787;
    defparam add_1980_3.INIT1 = 16'h7878;
    defparam add_1980_3.INJECT1_0 = "NO";
    defparam add_1980_3.INJECT1_1 = "NO";
    CCU2D add_1980_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(resetn_c), .B1(n21501), .C1(GND_net), .D1(GND_net), .COUT(n25115));   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam add_1980_1.INIT0 = 16'hF000;
    defparam add_1980_1.INIT1 = 16'h7777;
    defparam add_1980_1.INJECT1_0 = "NO";
    defparam add_1980_1.INJECT1_1 = "NO";
    FD1P3IX quad_set_valid_404 (.D(n29079), .SP(clk_enable_519), .CD(n29239), 
            .CK(clk), .Q(quad_set_valid)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=272, LSE_RLINE=293 */ ;   // c:/s_links/sources/quad_decoder.v(49[8] 63[4])
    defparam quad_set_valid_404.GSR = "DISABLED";
    LUT4 i16508_4_lut (.A(n2281[1]), .B(n29221), .C(n2281[3]), .D(n2281[2]), 
         .Z(n21446)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B (C+!(D))+!B !(C+!(D)))) */ ;
    defparam i16508_4_lut.init = 16'hc3c6;
    LUT4 i5163_4_lut (.A(n6171[0]), .B(quad_set[0]), .C(n5647), .D(n24), 
         .Z(n9956)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/s_links/sources/quad_decoder.v(124[18] 167[6])
    defparam i5163_4_lut.init = 16'hc0ca;
    
endmodule
//
// Verilog Description of module \stepper(DEV_ID=2,UART_ADDRESS_WIDTH=4) 
//

module \stepper(DEV_ID=2,UART_ADDRESS_WIDTH=4)  (clk_1MHz, clk_1MHz_enable_24, 
            n29239, mode_adj_134, clk, clk_enable_271, n29762, pin_io_out_29, 
            \quad_b[2] , pin_io_out_28, \quad_a[2] , spi_data_out_r_39__N_4496, 
            n47, digital_output_r, clk_enable_190, \spi_data_r[0] , 
            n29295, spi_data_out_r_39__N_4536, n19361, resetn_c, mode, 
            n29303, n22, GND_net, \spi_data_r[2] , \spi_data_r[1] , 
            n1, n8767, n29193, reset_r, clk_enable_306, n29070, 
            n1_adj_133, n29117, \spi_cmd[2] , n29212, n13413, quad_homing, 
            pin_io_out_24, n29233, n12714) /* synthesis syn_module_defined=1 */ ;
    input clk_1MHz;
    input clk_1MHz_enable_24;
    input n29239;
    output [2:0]mode_adj_134;
    input clk;
    input clk_enable_271;
    input n29762;
    input pin_io_out_29;
    output \quad_b[2] ;
    input pin_io_out_28;
    output \quad_a[2] ;
    output [39:0]spi_data_out_r_39__N_4496;
    input n47;
    output digital_output_r;
    input clk_enable_190;
    input \spi_data_r[0] ;
    output n29295;
    output spi_data_out_r_39__N_4536;
    output n19361;
    input resetn_c;
    input mode;
    input n29303;
    output n22;
    input GND_net;
    input \spi_data_r[2] ;
    input \spi_data_r[1] ;
    output n1;
    output n8767;
    output n29193;
    output reset_r;
    input clk_enable_306;
    input n29070;
    output n1_adj_133;
    input n29117;
    input \spi_cmd[2] ;
    input n29212;
    input n13413;
    input [1:0]quad_homing;
    input pin_io_out_24;
    input n29233;
    output n12714;
    
    wire clk_1MHz_derived_251 /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz_derived_251 */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire MA_Temp_N_4613 /* synthesis is_inv_clock=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire MA_Temp /* synthesis is_clock=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(57[5:12])
    wire [51:0]SLO;   // c:/s_links/sources/slot_cards/stepper.v(63[12:15])
    
    wire clk_1MHz_derived_251_enable_21;
    wire [51:0]SLO_buf;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    wire [11:0]Cnt_NSL;   // c:/s_links/sources/slot_cards/stepper.v(61[12:19])
    wire [11:0]n1290;
    wire [39:0]spi_data_out_r_39__N_4758;
    wire [7:0]Cnt;   // c:/s_links/sources/slot_cards/stepper.v(62[11:14])
    
    wire clk_1MHz_enable_73;
    wire [7:0]n199;
    
    wire n19429, n19509;
    wire [31:0]n153;
    
    wire n27334, n13366, n19457, n29297, n29257, spi_data_out_r_39__N_4829, 
        n29184, n11839, n29018, n29019, n29016, MA_Temp_N_4616, 
        n29017, clk_1MHz_enable_376, NSL, clk_1MHz_enable_101, NSL_N_4824, 
        n29139, n29296, n25004, n25003, n25002, n25001, n25000, 
        n24999, n24998, n24997, n24996, n24995, MA_Temp_N_4627, 
        clk_1MHz_derived_251_enable_46, n4;
    
    FD1P3AX SLO_i18 (.D(SLO[17]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i18.GSR = "DISABLED";
    FD1P3AX SLO_i17 (.D(SLO[16]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i17.GSR = "DISABLED";
    FD1P3AX SLO_i16 (.D(SLO[15]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i16.GSR = "DISABLED";
    FD1P3AX SLO_i15 (.D(SLO[14]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i15.GSR = "DISABLED";
    FD1P3AX SLO_i14 (.D(SLO[13]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i14.GSR = "DISABLED";
    FD1P3AX SLO_i13 (.D(SLO[12]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i13.GSR = "DISABLED";
    FD1P3AX SLO_i12 (.D(SLO[11]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i12.GSR = "DISABLED";
    FD1P3AX SLO_i11 (.D(SLO[10]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i11.GSR = "DISABLED";
    FD1P3AX SLO_i10 (.D(SLO[9]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i10.GSR = "DISABLED";
    FD1P3AX SLO_i9 (.D(SLO[8]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i9.GSR = "DISABLED";
    FD1P3AX SLO_i8 (.D(SLO[7]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i8.GSR = "DISABLED";
    FD1P3AX SLO_i7 (.D(SLO[6]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i7.GSR = "DISABLED";
    FD1P3AX SLO_i6 (.D(SLO[5]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i6.GSR = "DISABLED";
    FD1P3AX SLO_i5 (.D(SLO[4]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i5.GSR = "DISABLED";
    FD1P3AX SLO_i4 (.D(SLO[3]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i4.GSR = "DISABLED";
    FD1P3AX SLO_i3 (.D(SLO[2]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i3.GSR = "DISABLED";
    FD1P3AX SLO_i2 (.D(SLO[1]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i2.GSR = "DISABLED";
    FD1P3AX SLO_i1 (.D(SLO[0]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i1.GSR = "DISABLED";
    FD1S3AX SLO_buf_i46 (.D(SLO[45]), .CK(MA_Temp_N_4613), .Q(SLO_buf[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i46.GSR = "DISABLED";
    FD1S3AX SLO_buf_i45 (.D(SLO[44]), .CK(MA_Temp_N_4613), .Q(SLO_buf[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i45.GSR = "DISABLED";
    FD1S3AX SLO_buf_i44 (.D(SLO[43]), .CK(MA_Temp_N_4613), .Q(SLO_buf[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i44.GSR = "DISABLED";
    FD1S3AX SLO_buf_i43 (.D(SLO[42]), .CK(MA_Temp_N_4613), .Q(SLO_buf[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i43.GSR = "DISABLED";
    FD1S3AX SLO_buf_i42 (.D(SLO[41]), .CK(MA_Temp_N_4613), .Q(SLO_buf[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i42.GSR = "DISABLED";
    FD1S3AX SLO_buf_i41 (.D(SLO[40]), .CK(MA_Temp_N_4613), .Q(SLO_buf[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i41.GSR = "DISABLED";
    FD1S3AX SLO_buf_i40 (.D(SLO[39]), .CK(MA_Temp_N_4613), .Q(SLO_buf[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i40.GSR = "DISABLED";
    FD1S3AX SLO_buf_i39 (.D(SLO[38]), .CK(MA_Temp_N_4613), .Q(SLO_buf[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i39.GSR = "DISABLED";
    FD1S3AX SLO_buf_i38 (.D(SLO[37]), .CK(MA_Temp_N_4613), .Q(SLO_buf[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i38.GSR = "DISABLED";
    FD1S3AX SLO_buf_i37 (.D(SLO[36]), .CK(MA_Temp_N_4613), .Q(SLO_buf[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i37.GSR = "DISABLED";
    FD1S3AX SLO_buf_i36 (.D(SLO[35]), .CK(MA_Temp_N_4613), .Q(SLO_buf[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i36.GSR = "DISABLED";
    FD1S3AX SLO_buf_i35 (.D(SLO[34]), .CK(MA_Temp_N_4613), .Q(SLO_buf[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i35.GSR = "DISABLED";
    FD1S3AX SLO_buf_i34 (.D(SLO[33]), .CK(MA_Temp_N_4613), .Q(SLO_buf[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i34.GSR = "DISABLED";
    FD1S3AX SLO_buf_i33 (.D(SLO[32]), .CK(MA_Temp_N_4613), .Q(SLO_buf[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i33.GSR = "DISABLED";
    FD1S3AX SLO_buf_i32 (.D(SLO[31]), .CK(MA_Temp_N_4613), .Q(SLO_buf[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i32.GSR = "DISABLED";
    FD1S3AX SLO_buf_i31 (.D(SLO[30]), .CK(MA_Temp_N_4613), .Q(SLO_buf[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i31.GSR = "DISABLED";
    FD1S3AX SLO_buf_i30 (.D(SLO[29]), .CK(MA_Temp_N_4613), .Q(SLO_buf[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i30.GSR = "DISABLED";
    FD1S3AX SLO_buf_i29 (.D(SLO[28]), .CK(MA_Temp_N_4613), .Q(SLO_buf[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i29.GSR = "DISABLED";
    FD1S3AX SLO_buf_i28 (.D(SLO[27]), .CK(MA_Temp_N_4613), .Q(SLO_buf[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i28.GSR = "DISABLED";
    FD1S3AX SLO_buf_i27 (.D(SLO[26]), .CK(MA_Temp_N_4613), .Q(SLO_buf[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i27.GSR = "DISABLED";
    FD1S3AX SLO_buf_i26 (.D(SLO[25]), .CK(MA_Temp_N_4613), .Q(SLO_buf[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i26.GSR = "DISABLED";
    FD1S3AX SLO_buf_i25 (.D(SLO[24]), .CK(MA_Temp_N_4613), .Q(SLO_buf[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i25.GSR = "DISABLED";
    FD1S3AX SLO_buf_i24 (.D(SLO[23]), .CK(MA_Temp_N_4613), .Q(SLO_buf[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i24.GSR = "DISABLED";
    FD1S3AX SLO_buf_i23 (.D(SLO[22]), .CK(MA_Temp_N_4613), .Q(SLO_buf[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i23.GSR = "DISABLED";
    FD1S3AX SLO_buf_i22 (.D(SLO[21]), .CK(MA_Temp_N_4613), .Q(SLO_buf[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i22.GSR = "DISABLED";
    FD1S3AX SLO_buf_i21 (.D(SLO[20]), .CK(MA_Temp_N_4613), .Q(SLO_buf[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i21.GSR = "DISABLED";
    FD1S3AX SLO_buf_i20 (.D(SLO[19]), .CK(MA_Temp_N_4613), .Q(SLO_buf[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i20.GSR = "DISABLED";
    FD1S3AX SLO_buf_i19 (.D(SLO[18]), .CK(MA_Temp_N_4613), .Q(SLO_buf[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i19.GSR = "DISABLED";
    FD1S3AX SLO_buf_i18 (.D(SLO[17]), .CK(MA_Temp_N_4613), .Q(SLO_buf[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i18.GSR = "DISABLED";
    FD1S3AX SLO_buf_i17 (.D(SLO[16]), .CK(MA_Temp_N_4613), .Q(SLO_buf[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i17.GSR = "DISABLED";
    FD1S3AX SLO_buf_i16 (.D(SLO[15]), .CK(MA_Temp_N_4613), .Q(SLO_buf[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i16.GSR = "DISABLED";
    FD1S3AX SLO_buf_i15 (.D(SLO[14]), .CK(MA_Temp_N_4613), .Q(SLO_buf[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i15.GSR = "DISABLED";
    FD1S3AX SLO_buf_i14 (.D(SLO[13]), .CK(MA_Temp_N_4613), .Q(SLO_buf[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i14.GSR = "DISABLED";
    FD1S3AX SLO_buf_i13 (.D(SLO[12]), .CK(MA_Temp_N_4613), .Q(SLO_buf[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i13.GSR = "DISABLED";
    FD1S3AX SLO_buf_i12 (.D(SLO[11]), .CK(MA_Temp_N_4613), .Q(SLO_buf[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i12.GSR = "DISABLED";
    FD1S3AX SLO_buf_i11 (.D(SLO[10]), .CK(MA_Temp_N_4613), .Q(SLO_buf[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i11.GSR = "DISABLED";
    FD1S3AX SLO_buf_i10 (.D(SLO[9]), .CK(MA_Temp_N_4613), .Q(SLO_buf[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i10.GSR = "DISABLED";
    FD1S3AX SLO_buf_i9 (.D(SLO[8]), .CK(MA_Temp_N_4613), .Q(SLO_buf[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i9.GSR = "DISABLED";
    FD1S3AX SLO_buf_i8 (.D(SLO[7]), .CK(MA_Temp_N_4613), .Q(SLO_buf[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i8.GSR = "DISABLED";
    FD1S3AX SLO_buf_i7 (.D(SLO[6]), .CK(MA_Temp_N_4613), .Q(SLO_buf[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i7.GSR = "DISABLED";
    FD1S3AX SLO_buf_i6 (.D(SLO[5]), .CK(MA_Temp_N_4613), .Q(SLO_buf[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i6.GSR = "DISABLED";
    FD1S3AX SLO_buf_i5 (.D(SLO[4]), .CK(MA_Temp_N_4613), .Q(SLO_buf[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i5.GSR = "DISABLED";
    FD1S3AX SLO_buf_i4 (.D(SLO[3]), .CK(MA_Temp_N_4613), .Q(SLO_buf[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i4.GSR = "DISABLED";
    FD1S3AX SLO_buf_i3 (.D(SLO[2]), .CK(MA_Temp_N_4613), .Q(SLO_buf[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i3.GSR = "DISABLED";
    FD1S3AX SLO_buf_i2 (.D(SLO[1]), .CK(MA_Temp_N_4613), .Q(SLO_buf[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i2.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i11 (.D(n1290[11]), .SP(clk_1MHz_enable_24), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i11.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i10 (.D(n1290[10]), .SP(clk_1MHz_enable_24), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i10.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i9 (.D(n1290[9]), .SP(clk_1MHz_enable_24), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i9.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i8 (.D(n1290[8]), .SP(clk_1MHz_enable_24), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i8.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i7 (.D(n1290[7]), .SP(clk_1MHz_enable_24), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i7.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i6 (.D(n1290[6]), .SP(clk_1MHz_enable_24), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i6.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i5 (.D(n1290[5]), .SP(clk_1MHz_enable_24), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i5.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i4 (.D(n1290[4]), .SP(clk_1MHz_enable_24), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i4.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i3 (.D(n1290[3]), .SP(clk_1MHz_enable_24), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i3.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i2 (.D(n1290[2]), .SP(clk_1MHz_enable_24), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i2.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i1 (.D(n1290[1]), .SP(clk_1MHz_enable_24), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i1.GSR = "DISABLED";
    FD1P3IX mode__i0 (.D(n29762), .SP(clk_enable_271), .CD(n29239), .CK(clk), 
            .Q(mode_adj_134[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i0.GSR = "DISABLED";
    LUT4 Select_4098_i1_2_lut_4_lut (.A(mode_adj_134[0]), .B(mode_adj_134[1]), 
         .C(mode_adj_134[2]), .D(pin_io_out_29), .Z(\quad_b[2] )) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam Select_4098_i1_2_lut_4_lut.init = 16'h0400;
    LUT4 Select_4091_i1_2_lut_4_lut (.A(mode_adj_134[0]), .B(mode_adj_134[1]), 
         .C(mode_adj_134[2]), .D(pin_io_out_28), .Z(\quad_a[2] )) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam Select_4091_i1_2_lut_4_lut.init = 16'h0400;
    FD1P3IX Cnt_NSL__i0 (.D(n1290[0]), .SP(clk_1MHz_enable_24), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i0.GSR = "DISABLED";
    FD1S3AX SLO_buf_i1 (.D(SLO[0]), .CK(MA_Temp_N_4613), .Q(SLO_buf[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i1.GSR = "DISABLED";
    FD1P3AX SLO_i0 (.D(pin_io_out_28), .SP(clk_1MHz_derived_251_enable_21), 
            .CK(clk_1MHz_derived_251), .Q(SLO[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i0 (.D(spi_data_out_r_39__N_4758[0]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i0.GSR = "DISABLED";
    FD1P3IX Cnt__i0 (.D(n199[0]), .SP(clk_1MHz_enable_73), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i0.GSR = "DISABLED";
    FD1P3IX Cnt__i7 (.D(n199[7]), .SP(clk_1MHz_enable_73), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i7.GSR = "DISABLED";
    FD1P3IX Cnt__i6 (.D(n199[6]), .SP(clk_1MHz_enable_73), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i6.GSR = "DISABLED";
    FD1P3IX Cnt__i5 (.D(n199[5]), .SP(clk_1MHz_enable_73), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i5.GSR = "DISABLED";
    FD1P3IX Cnt__i4 (.D(n199[4]), .SP(clk_1MHz_enable_73), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i4.GSR = "DISABLED";
    FD1P3IX Cnt__i3 (.D(n199[3]), .SP(clk_1MHz_enable_73), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i3.GSR = "DISABLED";
    FD1P3IX Cnt__i2 (.D(n199[2]), .SP(clk_1MHz_enable_73), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i1 (.D(n199[1]), .SP(clk_1MHz_enable_73), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i1.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i39 (.D(SLO_buf[13]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i39.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i38 (.D(SLO_buf[12]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i38.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i37 (.D(SLO_buf[11]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i37.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i36 (.D(SLO_buf[10]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i36.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i35 (.D(spi_data_out_r_39__N_4758[35]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i35.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i34 (.D(spi_data_out_r_39__N_4758[34]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i34.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i33 (.D(spi_data_out_r_39__N_4758[33]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i33.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(spi_data_out_r_39__N_4758[32]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i31 (.D(SLO_buf[45]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i30 (.D(SLO_buf[44]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i29 (.D(SLO_buf[43]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i28 (.D(SLO_buf[42]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i27 (.D(SLO_buf[41]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i26 (.D(SLO_buf[40]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i25 (.D(SLO_buf[39]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i24 (.D(SLO_buf[38]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i23 (.D(SLO_buf[37]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i22 (.D(SLO_buf[36]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i21 (.D(SLO_buf[35]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i20 (.D(SLO_buf[34]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i19 (.D(SLO_buf[33]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i18 (.D(SLO_buf[32]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i17 (.D(SLO_buf[31]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i16 (.D(SLO_buf[30]), .CK(clk), .CD(n47), .Q(spi_data_out_r_39__N_4496[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(spi_data_out_r_39__N_4758[15]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(spi_data_out_r_39__N_4758[14]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(spi_data_out_r_39__N_4758[13]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(spi_data_out_r_39__N_4758[12]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(spi_data_out_r_39__N_4758[11]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(spi_data_out_r_39__N_4758[10]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(spi_data_out_r_39__N_4758[9]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(spi_data_out_r_39__N_4758[8]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(spi_data_out_r_39__N_4758[7]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(spi_data_out_r_39__N_4758[6]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(spi_data_out_r_39__N_4758[5]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(spi_data_out_r_39__N_4758[4]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(spi_data_out_r_39__N_4758[3]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(spi_data_out_r_39__N_4758[2]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(spi_data_out_r_39__N_4758[1]), .CK(clk), 
            .Q(spi_data_out_r_39__N_4496[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    LUT4 mux_149_i15_3_lut (.A(SLO_buf[28]), .B(SLO_buf[18]), .C(n47), 
         .Z(spi_data_out_r_39__N_4758[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i15_3_lut.init = 16'hcaca;
    LUT4 mux_149_i14_3_lut (.A(SLO_buf[27]), .B(SLO_buf[17]), .C(n47), 
         .Z(spi_data_out_r_39__N_4758[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i14_3_lut.init = 16'hcaca;
    LUT4 mux_149_i13_3_lut (.A(SLO_buf[26]), .B(SLO_buf[16]), .C(n47), 
         .Z(spi_data_out_r_39__N_4758[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i13_3_lut.init = 16'hcaca;
    LUT4 mux_149_i12_3_lut (.A(SLO_buf[25]), .B(SLO_buf[15]), .C(n47), 
         .Z(spi_data_out_r_39__N_4758[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i12_3_lut.init = 16'hcaca;
    LUT4 mux_149_i11_3_lut (.A(SLO_buf[24]), .B(SLO_buf[14]), .C(n47), 
         .Z(spi_data_out_r_39__N_4758[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i11_3_lut.init = 16'hcaca;
    LUT4 mux_149_i10_3_lut (.A(SLO_buf[23]), .B(SLO_buf[13]), .C(n47), 
         .Z(spi_data_out_r_39__N_4758[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i10_3_lut.init = 16'hcaca;
    LUT4 mux_149_i9_3_lut (.A(SLO_buf[22]), .B(SLO_buf[12]), .C(n47), 
         .Z(spi_data_out_r_39__N_4758[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i9_3_lut.init = 16'hcaca;
    LUT4 i13647_2_lut_3_lut (.A(n19429), .B(n19509), .C(n153[0]), .Z(n199[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13647_2_lut_3_lut.init = 16'h7070;
    LUT4 i13605_2_lut_3_lut (.A(n19429), .B(n19509), .C(n153[7]), .Z(n199[7])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13605_2_lut_3_lut.init = 16'h7070;
    LUT4 i13606_2_lut_3_lut (.A(n19429), .B(n19509), .C(n153[6]), .Z(n199[6])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13606_2_lut_3_lut.init = 16'h7070;
    LUT4 i13609_2_lut_3_lut (.A(n19429), .B(n19509), .C(n153[5]), .Z(n199[5])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13609_2_lut_3_lut.init = 16'h7070;
    LUT4 i13610_2_lut_3_lut (.A(n19429), .B(n19509), .C(n153[4]), .Z(n199[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13610_2_lut_3_lut.init = 16'h7070;
    LUT4 i13611_2_lut_3_lut (.A(n19429), .B(n19509), .C(n153[3]), .Z(n199[3])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13611_2_lut_3_lut.init = 16'h7070;
    LUT4 mux_149_i8_3_lut (.A(SLO_buf[21]), .B(SLO_buf[11]), .C(n47), 
         .Z(spi_data_out_r_39__N_4758[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i8_3_lut.init = 16'hcaca;
    LUT4 i13612_2_lut_3_lut (.A(n19429), .B(n19509), .C(n153[2]), .Z(n199[2])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13612_2_lut_3_lut.init = 16'h7070;
    LUT4 i13613_2_lut_3_lut (.A(n19429), .B(n19509), .C(n153[1]), .Z(n199[1])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13613_2_lut_3_lut.init = 16'h7070;
    LUT4 mux_149_i7_3_lut (.A(SLO_buf[20]), .B(SLO_buf[10]), .C(n47), 
         .Z(spi_data_out_r_39__N_4758[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i7_3_lut.init = 16'hcaca;
    LUT4 mux_149_i6_3_lut (.A(SLO_buf[19]), .B(SLO_buf[9]), .C(n47), .Z(spi_data_out_r_39__N_4758[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i6_3_lut.init = 16'hcaca;
    LUT4 mux_149_i5_3_lut (.A(SLO_buf[18]), .B(SLO_buf[8]), .C(n47), .Z(spi_data_out_r_39__N_4758[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i5_3_lut.init = 16'hcaca;
    LUT4 mux_149_i4_3_lut (.A(SLO_buf[17]), .B(SLO_buf[7]), .C(n47), .Z(spi_data_out_r_39__N_4758[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i4_3_lut.init = 16'hcaca;
    LUT4 mux_149_i3_3_lut (.A(SLO_buf[16]), .B(SLO_buf[6]), .C(n47), .Z(spi_data_out_r_39__N_4758[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i3_3_lut.init = 16'hcaca;
    LUT4 mux_149_i2_3_lut (.A(SLO_buf[15]), .B(SLO_buf[5]), .C(n47), .Z(spi_data_out_r_39__N_4758[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i2_3_lut.init = 16'hcaca;
    FD1P3IX digital_output_r_481 (.D(\spi_data_r[0] ), .SP(clk_enable_190), 
            .CD(n29239), .CK(clk), .Q(digital_output_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam digital_output_r_481.GSR = "DISABLED";
    LUT4 i2_4_lut (.A(n27334), .B(Cnt[5]), .C(n13366), .D(n19457), .Z(n19429)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i2_4_lut.init = 16'hfefa;
    LUT4 i3_4_lut (.A(n19457), .B(Cnt[5]), .C(n29295), .D(n27334), .Z(n19509)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(Cnt[6]), .B(Cnt[7]), .Z(n27334)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i14517_4_lut (.A(Cnt[0]), .B(Cnt[4]), .C(n29297), .D(Cnt[1]), 
         .Z(n19457)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i14517_4_lut.init = 16'hc8c0;
    LUT4 i14322_2_lut_rep_529 (.A(Cnt[4]), .B(Cnt[1]), .Z(n29257)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14322_2_lut_rep_529.init = 16'h8888;
    FD1S3IX i159_483 (.D(spi_data_out_r_39__N_4829), .CK(clk), .CD(n29239), 
            .Q(spi_data_out_r_39__N_4536)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam i159_483.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(n29184), .D(Cnt[5]), 
         .Z(n11839)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff7;
    LUT4 n19429_bdd_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(Cnt[5]), .D(MA_Temp), 
         .Z(n29018)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;
    defparam n19429_bdd_3_lut_4_lut.init = 16'hf708;
    LUT4 n29019_bdd_3_lut (.A(n29019), .B(n29016), .C(n29184), .Z(MA_Temp_N_4616)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n29019_bdd_3_lut.init = 16'hcaca;
    LUT4 n19429_bdd_3_lut_23138 (.A(n19429), .B(n19509), .C(MA_Temp), 
         .Z(n29016)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam n19429_bdd_3_lut_23138.init = 16'h7070;
    LUT4 n19429_bdd_4_lut_23345 (.A(n19429), .B(n29257), .C(MA_Temp), 
         .D(Cnt[5]), .Z(n29017)) /* synthesis lut_function=(!(A+(B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam n19429_bdd_4_lut_23345.init = 16'h1450;
    LUT4 i22827_2_lut_rep_437 (.A(n19361), .B(resetn_c), .Z(clk_1MHz_enable_73)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i22827_2_lut_rep_437.init = 16'hbbbb;
    LUT4 i22868_2_lut_2_lut_3_lut_4_lut (.A(n19361), .B(resetn_c), .C(n19509), 
         .D(n19429), .Z(clk_1MHz_enable_376)) /* synthesis lut_function=(!(A (C (D))+!A (B+(C (D))))) */ ;
    defparam i22868_2_lut_2_lut_3_lut_4_lut.init = 16'h0bbb;
    FD1P3AX NSL_476 (.D(NSL_N_4824), .SP(clk_1MHz_enable_101), .CK(clk_1MHz), 
            .Q(NSL)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam NSL_476.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_411_4_lut (.A(n29297), .B(Cnt[0]), .C(n27334), .D(Cnt[5]), 
         .Z(n29139)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_rep_411_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_4_lut (.A(mode_adj_134[2]), .B(n29296), .C(mode), .D(n29303), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    CCU2D add_551_13 (.A0(Cnt_NSL[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25004), 
          .S0(n1290[11]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_13.INIT0 = 16'h5aaa;
    defparam add_551_13.INIT1 = 16'h0000;
    defparam add_551_13.INJECT1_0 = "NO";
    defparam add_551_13.INJECT1_1 = "NO";
    CCU2D add_551_11 (.A0(Cnt_NSL[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25003), .COUT(n25004), .S0(n1290[9]), .S1(n1290[10]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_11.INIT0 = 16'h5aaa;
    defparam add_551_11.INIT1 = 16'h5aaa;
    defparam add_551_11.INJECT1_0 = "NO";
    defparam add_551_11.INJECT1_1 = "NO";
    CCU2D add_551_9 (.A0(Cnt_NSL[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25002), .COUT(n25003), .S0(n1290[7]), .S1(n1290[8]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_9.INIT0 = 16'h5aaa;
    defparam add_551_9.INIT1 = 16'h5aaa;
    defparam add_551_9.INJECT1_0 = "NO";
    defparam add_551_9.INJECT1_1 = "NO";
    CCU2D add_551_7 (.A0(Cnt_NSL[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25001), .COUT(n25002), .S0(n1290[5]), .S1(n1290[6]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_7.INIT0 = 16'h5aaa;
    defparam add_551_7.INIT1 = 16'h5aaa;
    defparam add_551_7.INJECT1_0 = "NO";
    defparam add_551_7.INJECT1_1 = "NO";
    CCU2D add_551_5 (.A0(Cnt_NSL[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25000), .COUT(n25001), .S0(n1290[3]), .S1(n1290[4]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_5.INIT0 = 16'h5aaa;
    defparam add_551_5.INIT1 = 16'h5aaa;
    defparam add_551_5.INJECT1_0 = "NO";
    defparam add_551_5.INJECT1_1 = "NO";
    CCU2D add_551_3 (.A0(Cnt_NSL[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24999), .COUT(n25000), .S0(n1290[1]), .S1(n1290[2]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_3.INIT0 = 16'h5aaa;
    defparam add_551_3.INIT1 = 16'h5aaa;
    defparam add_551_3.INJECT1_0 = "NO";
    defparam add_551_3.INJECT1_1 = "NO";
    FD1P3IX mode__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_271), .CD(n29239), 
            .CK(clk), .Q(mode_adj_134[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i2.GSR = "DISABLED";
    FD1P3IX mode__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_271), .CD(n29239), 
            .CK(clk), .Q(mode_adj_134[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i1.GSR = "DISABLED";
    CCU2D add_551_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24999), .S1(n1290[0]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_1.INIT0 = 16'hF000;
    defparam add_551_1.INIT1 = 16'h5555;
    defparam add_551_1.INJECT1_0 = "NO";
    defparam add_551_1.INJECT1_1 = "NO";
    CCU2D add_552_9 (.A0(Cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24998), 
          .S0(n153[7]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_9.INIT0 = 16'h5aaa;
    defparam add_552_9.INIT1 = 16'h0000;
    defparam add_552_9.INJECT1_0 = "NO";
    defparam add_552_9.INJECT1_1 = "NO";
    LUT4 mux_149_i1_3_lut (.A(SLO_buf[14]), .B(SLO_buf[4]), .C(n47), .Z(spi_data_out_r_39__N_4758[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i1_3_lut.init = 16'hcaca;
    CCU2D add_552_7 (.A0(Cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24997), 
          .COUT(n24998), .S0(n153[5]), .S1(n153[6]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_7.INIT0 = 16'h5aaa;
    defparam add_552_7.INIT1 = 16'h5aaa;
    defparam add_552_7.INJECT1_0 = "NO";
    defparam add_552_7.INJECT1_1 = "NO";
    CCU2D add_552_5 (.A0(Cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24996), 
          .COUT(n24997), .S0(n153[3]), .S1(n153[4]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_5.INIT0 = 16'h5aaa;
    defparam add_552_5.INIT1 = 16'h5aaa;
    defparam add_552_5.INJECT1_0 = "NO";
    defparam add_552_5.INJECT1_1 = "NO";
    CCU2D add_552_3 (.A0(Cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24995), 
          .COUT(n24996), .S0(n153[1]), .S1(n153[2]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_3.INIT0 = 16'h5aaa;
    defparam add_552_3.INIT1 = 16'h5aaa;
    defparam add_552_3.INJECT1_0 = "NO";
    defparam add_552_3.INJECT1_1 = "NO";
    CCU2D add_552_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24995), 
          .S1(n153[0]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_1.INIT0 = 16'hF000;
    defparam add_552_1.INIT1 = 16'h5555;
    defparam add_552_1.INJECT1_0 = "NO";
    defparam add_552_1.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_567 (.A(mode_adj_134[2]), .B(mode_adj_134[0]), .C(mode_adj_134[1]), 
         .Z(n29295)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i2_3_lut_rep_567.init = 16'hf7f7;
    LUT4 Select_3966_i1_2_lut_4_lut (.A(mode_adj_134[2]), .B(mode_adj_134[0]), 
         .C(mode_adj_134[1]), .D(NSL), .Z(n1)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam Select_3966_i1_2_lut_4_lut.init = 16'h0800;
    LUT4 i22723_2_lut_2_lut_4_lut (.A(mode_adj_134[2]), .B(mode_adj_134[0]), 
         .C(mode_adj_134[1]), .D(n29303), .Z(n8767)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i22723_2_lut_2_lut_4_lut.init = 16'h00f7;
    LUT4 equal_115_i6_1_lut_3_lut (.A(mode_adj_134[2]), .B(mode_adj_134[0]), 
         .C(mode_adj_134[1]), .Z(MA_Temp_N_4627)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam equal_115_i6_1_lut_3_lut.init = 16'h0808;
    LUT4 i4788_2_lut_4_lut (.A(mode_adj_134[2]), .B(mode_adj_134[0]), .C(mode_adj_134[1]), 
         .D(clk_1MHz_derived_251_enable_46), .Z(clk_1MHz_derived_251_enable_21)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (D)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i4788_2_lut_4_lut.init = 16'hff08;
    LUT4 i1_2_lut_rep_568 (.A(mode_adj_134[1]), .B(mode_adj_134[0]), .Z(n29296)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_rep_568.init = 16'heeee;
    LUT4 i1_2_lut_rep_465_3_lut (.A(mode_adj_134[1]), .B(mode_adj_134[0]), 
         .C(mode_adj_134[2]), .Z(n29193)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_rep_465_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut (.A(mode_adj_134[1]), .B(mode_adj_134[0]), .C(mode_adj_134[2]), 
         .Z(n13366)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_569 (.A(Cnt[2]), .B(Cnt[3]), .Z(n29297)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_rep_569.init = 16'heeee;
    LUT4 i2_3_lut_rep_456_4_lut (.A(Cnt[2]), .B(Cnt[3]), .C(n27334), .D(Cnt[0]), 
         .Z(n29184)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i2_3_lut_rep_456_4_lut.init = 16'hfffe;
    FD1P3IX SLO_i45 (.D(SLO[44]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i45.GSR = "DISABLED";
    FD1P3IX reset_r_480 (.D(n29070), .SP(clk_enable_306), .CD(n29239), 
            .CK(clk), .Q(reset_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam reset_r_480.GSR = "DISABLED";
    FD1P3AX SLO_i19 (.D(SLO[18]), .SP(clk_1MHz_derived_251_enable_21), .CK(clk_1MHz_derived_251), 
            .Q(SLO[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i19.GSR = "DISABLED";
    FD1P3IX SLO_i44 (.D(SLO[43]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i44.GSR = "DISABLED";
    FD1P3IX SLO_i43 (.D(SLO[42]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i43.GSR = "DISABLED";
    FD1P3IX SLO_i42 (.D(SLO[41]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i42.GSR = "DISABLED";
    FD1P3IX SLO_i41 (.D(SLO[40]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i41.GSR = "DISABLED";
    FD1P3IX SLO_i40 (.D(SLO[39]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i40.GSR = "DISABLED";
    FD1P3IX SLO_i39 (.D(SLO[38]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i39.GSR = "DISABLED";
    FD1P3IX SLO_i38 (.D(SLO[37]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i38.GSR = "DISABLED";
    FD1P3IX SLO_i37 (.D(SLO[36]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i37.GSR = "DISABLED";
    FD1P3IX SLO_i36 (.D(SLO[35]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i36.GSR = "DISABLED";
    FD1P3IX SLO_i35 (.D(SLO[34]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i35.GSR = "DISABLED";
    FD1P3IX SLO_i34 (.D(SLO[33]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i34.GSR = "DISABLED";
    FD1P3IX SLO_i33 (.D(SLO[32]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i33.GSR = "DISABLED";
    FD1P3IX SLO_i32 (.D(SLO[31]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i32.GSR = "DISABLED";
    FD1P3IX SLO_i31 (.D(SLO[30]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i31.GSR = "DISABLED";
    FD1P3IX SLO_i30 (.D(SLO[29]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i30.GSR = "DISABLED";
    FD1P3IX SLO_i29 (.D(SLO[28]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i29.GSR = "DISABLED";
    FD1P3IX SLO_i28 (.D(SLO[27]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i28.GSR = "DISABLED";
    FD1P3IX SLO_i27 (.D(SLO[26]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i27.GSR = "DISABLED";
    FD1P3IX SLO_i26 (.D(SLO[25]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i26.GSR = "DISABLED";
    FD1P3IX SLO_i25 (.D(SLO[24]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i25.GSR = "DISABLED";
    FD1P3IX SLO_i24 (.D(SLO[23]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i24.GSR = "DISABLED";
    FD1P3IX SLO_i23 (.D(SLO[22]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i23.GSR = "DISABLED";
    FD1P3IX SLO_i22 (.D(SLO[21]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i22.GSR = "DISABLED";
    FD1P3IX SLO_i21 (.D(SLO[20]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i21.GSR = "DISABLED";
    FD1P3IX SLO_i20 (.D(SLO[19]), .SP(clk_1MHz_derived_251_enable_46), .CD(MA_Temp_N_4627), 
            .CK(clk_1MHz_derived_251), .Q(SLO[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i20.GSR = "DISABLED";
    LUT4 mux_149_i33_3_lut (.A(SLO_buf[6]), .B(SLO_buf[0]), .C(n47), .Z(spi_data_out_r_39__N_4758[32])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i33_3_lut.init = 16'hcaca;
    FD1P3IX MA_Temp_474 (.D(MA_Temp_N_4616), .SP(clk_1MHz_enable_376), .CD(n29239), 
            .CK(clk_1MHz), .Q(MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam MA_Temp_474.GSR = "DISABLED";
    LUT4 i22638_2_lut_rep_586 (.A(MA_Temp), .B(clk_1MHz), .Z(clk_1MHz_derived_251)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[13:34])
    defparam i22638_2_lut_rep_586.init = 16'h7777;
    LUT4 Select_3963_i1_2_lut_3_lut (.A(MA_Temp), .B(clk_1MHz), .C(mode_adj_134[2]), 
         .Z(n1_adj_133)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[13:34])
    defparam Select_3963_i1_2_lut_3_lut.init = 16'h7070;
    LUT4 i117_4_lut (.A(n29139), .B(n13366), .C(Cnt[4]), .D(Cnt[1]), 
         .Z(clk_1MHz_derived_251_enable_46)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(132[15:49])
    defparam i117_4_lut.init = 16'h3332;
    LUT4 i22641_4_lut (.A(n29117), .B(\spi_cmd[2] ), .C(n29212), .D(n13413), 
         .Z(spi_data_out_r_39__N_4829)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;
    defparam i22641_4_lut.init = 16'h0444;
    LUT4 i3_4_lut_adj_480 (.A(quad_homing[0]), .B(quad_homing[1]), .C(pin_io_out_24), 
         .D(n29233), .Z(n12714)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(75[8:17])
    defparam i3_4_lut_adj_480.init = 16'h0020;
    LUT4 i14347_3_lut (.A(n19509), .B(resetn_c), .C(n19361), .Z(clk_1MHz_enable_101)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B))) */ ;
    defparam i14347_3_lut.init = 16'h4c4c;
    LUT4 i22635_4_lut (.A(NSL), .B(n19361), .C(n19509), .D(n11839), 
         .Z(NSL_N_4824)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C+(D))))) */ ;
    defparam i22635_4_lut.init = 16'h3b37;
    LUT4 i2_4_lut_adj_481 (.A(Cnt_NSL[11]), .B(Cnt_NSL[9]), .C(Cnt_NSL[10]), 
         .D(n4), .Z(n19361)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_481.init = 16'ha080;
    LUT4 i1_2_lut_adj_482 (.A(Cnt_NSL[7]), .B(Cnt_NSL[8]), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_482.init = 16'heeee;
    PFUMX i23139 (.BLUT(n29018), .ALUT(n29017), .C0(n19509), .Z(n29019));
    LUT4 mux_149_i36_3_lut (.A(SLO_buf[9]), .B(SLO_buf[3]), .C(n47), .Z(spi_data_out_r_39__N_4758[35])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i36_3_lut.init = 16'hcaca;
    LUT4 mux_149_i35_3_lut (.A(SLO_buf[8]), .B(SLO_buf[2]), .C(n47), .Z(spi_data_out_r_39__N_4758[34])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i35_3_lut.init = 16'hcaca;
    LUT4 mux_149_i34_3_lut (.A(SLO_buf[7]), .B(SLO_buf[1]), .C(n47), .Z(spi_data_out_r_39__N_4758[33])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i34_3_lut.init = 16'hcaca;
    INV i23371 (.A(MA_Temp), .Z(MA_Temp_N_4613));
    LUT4 mux_149_i16_3_lut (.A(SLO_buf[29]), .B(SLO_buf[19]), .C(n47), 
         .Z(spi_data_out_r_39__N_4758[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[11] 208[5])
    defparam mux_149_i16_3_lut.init = 16'hcaca;
    
endmodule
//
// Verilog Description of module \stepper(UART_ADDRESS_WIDTH=4) 
//

module \stepper(UART_ADDRESS_WIDTH=4)  (\spi_cmd[0] , n29108, \SLO_buf[4] , 
            \SLO_buf[14] , \spi_data_out_r_39__N_5775[0] , \SLO_buf[3] , 
            \SLO_buf[9] , \spi_data_out_r_39__N_5775[35] , \SLO_buf[2] , 
            \SLO_buf[8] , \spi_data_out_r_39__N_5775[34] , \SLO_buf[1] , 
            \SLO_buf[7] , \spi_data_out_r_39__N_5775[33] , n29087, \SLO_buf[16] , 
            \SLO_buf[26] , \spi_data_out_r_39__N_6114[12] , \SLO_buf[0] , 
            \SLO_buf[6] , \spi_data_out_r_39__N_5775[32] , \SLO_buf[19] , 
            \SLO_buf[29] , \spi_data_out_r_39__N_5775[15] , \SLO_buf[18] , 
            \SLO_buf[28] , \spi_data_out_r_39__N_5775[14] , \SLO_buf[17] , 
            \SLO_buf[27] , \spi_data_out_r_39__N_5775[13] , \SLO_buf[16]_adj_11 , 
            \SLO_buf[26]_adj_12 , \spi_data_out_r_39__N_5775[12] , \SLO_buf[15] , 
            \SLO_buf[25] , \spi_data_out_r_39__N_5775[11] , \SLO_buf[24] , 
            \spi_data_out_r_39__N_5775[10] , \SLO_buf[13] , \SLO_buf[23] , 
            \spi_data_out_r_39__N_5775[9] , \SLO_buf[12] , \SLO_buf[22] , 
            \spi_data_out_r_39__N_5775[8] , \SLO_buf[11] , \SLO_buf[21] , 
            \spi_data_out_r_39__N_5775[7] , \SLO_buf[10] , \SLO_buf[20] , 
            \spi_data_out_r_39__N_5775[6] , \spi_data_out_r_39__N_5775[5] , 
            \spi_data_out_r_39__N_5775[4] , \spi_data_out_r_39__N_5775[3] , 
            \spi_data_out_r_39__N_5775[2] , pin_io_out_8, spi_data_out_r_39__N_3818, 
            clk, \SLO_buf[5] , \spi_data_out_r_39__N_5775[1] , mode_adj_132, 
            clk_1MHz, n29239, pin_io_out_9, \quad_b[0] , \quad_a[0] , 
            n29201, clk_1MHz_enable_55, clk_enable_402, n29762, n29185, 
            \spi_addr[1] , n29761, \spi_addr[2] , \spi_cmd[2] , n13489, 
            n29178, digital_output_r, clk_enable_173, \spi_data_r[0] , 
            spi_data_out_r_39__N_3858, \SLO_buf[4]_adj_13 , \SLO_buf[14]_adj_14 , 
            \spi_data_out_r_39__N_6114[0] , \SLO_buf[3]_adj_15 , \SLO_buf[9]_adj_16 , 
            \spi_data_out_r_39__N_6114[35] , resetn_c, n19337, \SLO_buf[15]_adj_17 , 
            \SLO_buf[25]_adj_18 , \spi_data_out_r_39__N_6114[11] , \SLO_buf[24]_adj_19 , 
            \spi_data_out_r_39__N_6114[10] , \SLO_buf[13]_adj_20 , \SLO_buf[23]_adj_21 , 
            \spi_data_out_r_39__N_6114[9] , \SLO_buf[4]_adj_22 , \SLO_buf[14]_adj_23 , 
            \spi_data_out_r_39__N_5436[0] , \SLO_buf[3]_adj_24 , \SLO_buf[9]_adj_25 , 
            \spi_data_out_r_39__N_5436[35] , \SLO_buf[2]_adj_26 , \SLO_buf[8]_adj_27 , 
            \spi_data_out_r_39__N_6114[34] , \SLO_buf[2]_adj_28 , \SLO_buf[8]_adj_29 , 
            \spi_data_out_r_39__N_5436[34] , \SLO_buf[1]_adj_30 , \SLO_buf[7]_adj_31 , 
            \spi_data_out_r_39__N_5436[33] , \SLO_buf[0]_adj_32 , \SLO_buf[6]_adj_33 , 
            \spi_data_out_r_39__N_5436[32] , \SLO_buf[12]_adj_34 , \SLO_buf[22]_adj_35 , 
            \spi_data_out_r_39__N_6114[8] , \SLO_buf[19]_adj_36 , \SLO_buf[29]_adj_37 , 
            \spi_data_out_r_39__N_5436[15] , \SLO_buf[18]_adj_38 , \SLO_buf[28]_adj_39 , 
            \spi_data_out_r_39__N_5436[14] , \SLO_buf[11]_adj_40 , \SLO_buf[21]_adj_41 , 
            \spi_data_out_r_39__N_6114[7] , \SLO_buf[10]_adj_42 , \SLO_buf[20]_adj_43 , 
            \spi_data_out_r_39__N_6114[6] , \SLO_buf[17]_adj_44 , \SLO_buf[27]_adj_45 , 
            \spi_data_out_r_39__N_5436[13] , \SLO_buf[16]_adj_46 , \SLO_buf[26]_adj_47 , 
            \spi_data_out_r_39__N_5436[12] , \SLO_buf[15]_adj_48 , \SLO_buf[25]_adj_49 , 
            \spi_data_out_r_39__N_5436[11] , \SLO_buf[1]_adj_50 , \SLO_buf[7]_adj_51 , 
            \spi_data_out_r_39__N_6114[33] , \SLO_buf[24]_adj_52 , \spi_data_out_r_39__N_5436[10] , 
            \SLO_buf[13]_adj_53 , \SLO_buf[23]_adj_54 , \spi_data_out_r_39__N_5436[9] , 
            n1, \SLO_buf[0]_adj_55 , \SLO_buf[6]_adj_56 , \spi_data_out_r_39__N_6114[32] , 
            n29309, n8823, n29216, n29205, \spi_addr_r[1] , n29214, 
            n29134, \SLO_buf[12]_adj_57 , \SLO_buf[22]_adj_58 , \spi_data_out_r_39__N_5436[8] , 
            \SLO_buf[11]_adj_59 , \SLO_buf[21]_adj_60 , \spi_data_out_r_39__N_5436[7] , 
            \SLO_buf[10]_adj_61 , \SLO_buf[20]_adj_62 , \spi_data_out_r_39__N_5436[6] , 
            \spi_data_out_r_39__N_5436[5] , \spi_data_out_r_39__N_5436[4] , 
            \spi_data_out_r_39__N_5436[3] , \spi_data_out_r_39__N_5436[2] , 
            \SLO_buf[19]_adj_63 , \SLO_buf[29]_adj_64 , \spi_data_out_r_39__N_6114[15] , 
            n1_adj_65, \cs_decoded[0] , n8824, \SLO_buf[5]_adj_66 , 
            \spi_data_out_r_39__N_5436[1] , \spi_data_out_r_39__N_6114[5] , 
            n18550, \SLO_buf[18]_adj_67 , \spi_data_out_r_39__N_6114[4] , 
            GND_net, n29310, \SLO_buf[4]_adj_68 , \SLO_buf[14]_adj_69 , 
            \spi_data_out_r_39__N_5097[0] , \SLO_buf[3]_adj_70 , \SLO_buf[9]_adj_71 , 
            \spi_data_out_r_39__N_5097[35] , \SLO_buf[2]_adj_72 , \SLO_buf[8]_adj_73 , 
            \spi_data_out_r_39__N_5097[34] , \SLO_buf[17]_adj_74 , \spi_data_out_r_39__N_6114[3] , 
            \spi_data_out_r_39__N_6114[2] , \SLO_buf[28]_adj_75 , \spi_data_out_r_39__N_6114[14] , 
            mode, n31, n22, \SLO_buf[1]_adj_76 , \SLO_buf[7]_adj_77 , 
            \spi_data_out_r_39__N_5097[33] , \SLO_buf[0]_adj_78 , \SLO_buf[6]_adj_79 , 
            \spi_data_out_r_39__N_5097[32] , \SLO_buf[5]_adj_80 , \spi_data_out_r_39__N_6114[1] , 
            \SLO_buf[19]_adj_81 , \SLO_buf[29]_adj_82 , \spi_data_out_r_39__N_5097[15] , 
            \SLO_buf[18]_adj_83 , \SLO_buf[28]_adj_84 , \spi_data_out_r_39__N_5097[14] , 
            \SLO_buf[17]_adj_85 , \SLO_buf[27]_adj_86 , \spi_data_out_r_39__N_5097[13] , 
            \SLO_buf[16]_adj_87 , \SLO_buf[26]_adj_88 , \spi_data_out_r_39__N_5097[12] , 
            \SLO_buf[15]_adj_89 , \SLO_buf[25]_adj_90 , \spi_data_out_r_39__N_5097[11] , 
            \SLO_buf[24]_adj_91 , \spi_data_out_r_39__N_5097[10] , \SLO_buf[13]_adj_92 , 
            \SLO_buf[23]_adj_93 , \spi_data_out_r_39__N_5097[9] , \SLO_buf[12]_adj_94 , 
            \SLO_buf[22]_adj_95 , \spi_data_out_r_39__N_5097[8] , \SLO_buf[11]_adj_96 , 
            \SLO_buf[21]_adj_97 , \spi_data_out_r_39__N_5097[7] , \SLO_buf[10]_adj_98 , 
            \SLO_buf[20]_adj_99 , \spi_data_out_r_39__N_5097[6] , \spi_cmd_r[1] , 
            \spi_addr_r[0] , n29287, \spi_cmd_r[0] , n29311, n27286, 
            \SLO_buf[27]_adj_100 , \spi_data_out_r_39__N_6114[13] , \spi_data_out_r_39__N_5097[5] , 
            \spi_data_out_r_39__N_5097[4] , \spi_data_out_r_39__N_5097[3] , 
            \spi_data_out_r_39__N_5097[2] , \SLO_buf[5]_adj_101 , \spi_data_out_r_39__N_5097[1] , 
            \SLO_buf[3]_adj_102 , \SLO_buf[9]_adj_103 , \spi_data_out_r_39__N_4419[35] , 
            \SLO_buf[2]_adj_104 , \SLO_buf[8]_adj_105 , \spi_data_out_r_39__N_4419[34] , 
            \SLO_buf[1]_adj_106 , \SLO_buf[7]_adj_107 , \spi_data_out_r_39__N_4419[33] , 
            \SLO_buf[0]_adj_108 , \SLO_buf[6]_adj_109 , \spi_data_out_r_39__N_4419[32] , 
            \SLO_buf[19]_adj_110 , \SLO_buf[29]_adj_111 , \spi_data_out_r_39__N_4419[15] , 
            \SLO_buf[18]_adj_112 , \SLO_buf[28]_adj_113 , \spi_data_out_r_39__N_4419[14] , 
            \SLO_buf[17]_adj_114 , \SLO_buf[27]_adj_115 , \spi_data_out_r_39__N_4419[13] , 
            \SLO_buf[16]_adj_116 , \SLO_buf[26]_adj_117 , \spi_data_out_r_39__N_4419[12] , 
            \SLO_buf[15]_adj_118 , \SLO_buf[25]_adj_119 , \spi_data_out_r_39__N_4419[11] , 
            \SLO_buf[14]_adj_120 , \SLO_buf[24]_adj_121 , \spi_data_out_r_39__N_4419[10] , 
            \SLO_buf[13]_adj_122 , \SLO_buf[23]_adj_123 , \spi_data_out_r_39__N_4419[9] , 
            \SLO_buf[12]_adj_124 , \SLO_buf[22]_adj_125 , \spi_data_out_r_39__N_4419[8] , 
            \SLO_buf[11]_adj_126 , \SLO_buf[21]_adj_127 , \spi_data_out_r_39__N_4419[7] , 
            \SLO_buf[10]_adj_128 , \SLO_buf[20]_adj_129 , \spi_data_out_r_39__N_4419[6] , 
            \spi_data_out_r_39__N_4419[5] , \spi_data_out_r_39__N_4419[4] , 
            \spi_data_out_r_39__N_4419[3] , \spi_data_out_r_39__N_4419[2] , 
            \SLO_buf[5]_adj_130 , \spi_data_out_r_39__N_4419[1] , \SLO_buf[4]_adj_131 , 
            \spi_data_out_r_39__N_4419[0] , \spi_data_r[1] , \spi_data_r[2] , 
            reset_r, clk_enable_506, n29106, n29117, n29076, n29115, 
            spi_data_out_r_39__N_4490, n29093, n29094, \spi_addr[0] , 
            n29126, clear_intrpt_N_2710, \spi_cmd[1] , n29141, n26933, 
            n29212, n47, clear_intrpt_N_2639, spi_data_out_r_39__N_5507, 
            n29091, n29098, n29099) /* synthesis syn_module_defined=1 */ ;
    input \spi_cmd[0] ;
    output n29108;
    input \SLO_buf[4] ;
    input \SLO_buf[14] ;
    output \spi_data_out_r_39__N_5775[0] ;
    input \SLO_buf[3] ;
    input \SLO_buf[9] ;
    output \spi_data_out_r_39__N_5775[35] ;
    input \SLO_buf[2] ;
    input \SLO_buf[8] ;
    output \spi_data_out_r_39__N_5775[34] ;
    input \SLO_buf[1] ;
    input \SLO_buf[7] ;
    output \spi_data_out_r_39__N_5775[33] ;
    output n29087;
    input \SLO_buf[16] ;
    input \SLO_buf[26] ;
    output \spi_data_out_r_39__N_6114[12] ;
    input \SLO_buf[0] ;
    input \SLO_buf[6] ;
    output \spi_data_out_r_39__N_5775[32] ;
    input \SLO_buf[19] ;
    input \SLO_buf[29] ;
    output \spi_data_out_r_39__N_5775[15] ;
    input \SLO_buf[18] ;
    input \SLO_buf[28] ;
    output \spi_data_out_r_39__N_5775[14] ;
    input \SLO_buf[17] ;
    input \SLO_buf[27] ;
    output \spi_data_out_r_39__N_5775[13] ;
    input \SLO_buf[16]_adj_11 ;
    input \SLO_buf[26]_adj_12 ;
    output \spi_data_out_r_39__N_5775[12] ;
    input \SLO_buf[15] ;
    input \SLO_buf[25] ;
    output \spi_data_out_r_39__N_5775[11] ;
    input \SLO_buf[24] ;
    output \spi_data_out_r_39__N_5775[10] ;
    input \SLO_buf[13] ;
    input \SLO_buf[23] ;
    output \spi_data_out_r_39__N_5775[9] ;
    input \SLO_buf[12] ;
    input \SLO_buf[22] ;
    output \spi_data_out_r_39__N_5775[8] ;
    input \SLO_buf[11] ;
    input \SLO_buf[21] ;
    output \spi_data_out_r_39__N_5775[7] ;
    input \SLO_buf[10] ;
    input \SLO_buf[20] ;
    output \spi_data_out_r_39__N_5775[6] ;
    output \spi_data_out_r_39__N_5775[5] ;
    output \spi_data_out_r_39__N_5775[4] ;
    output \spi_data_out_r_39__N_5775[3] ;
    output \spi_data_out_r_39__N_5775[2] ;
    input pin_io_out_8;
    output [39:0]spi_data_out_r_39__N_3818;
    input clk;
    input \SLO_buf[5] ;
    output \spi_data_out_r_39__N_5775[1] ;
    output [2:0]mode_adj_132;
    input clk_1MHz;
    input n29239;
    input pin_io_out_9;
    output \quad_b[0] ;
    output \quad_a[0] ;
    output n29201;
    input clk_1MHz_enable_55;
    input clk_enable_402;
    input n29762;
    output n29185;
    input \spi_addr[1] ;
    input n29761;
    input \spi_addr[2] ;
    input \spi_cmd[2] ;
    output n13489;
    output n29178;
    output digital_output_r;
    input clk_enable_173;
    input \spi_data_r[0] ;
    output spi_data_out_r_39__N_3858;
    input \SLO_buf[4]_adj_13 ;
    input \SLO_buf[14]_adj_14 ;
    output \spi_data_out_r_39__N_6114[0] ;
    input \SLO_buf[3]_adj_15 ;
    input \SLO_buf[9]_adj_16 ;
    output \spi_data_out_r_39__N_6114[35] ;
    input resetn_c;
    output n19337;
    input \SLO_buf[15]_adj_17 ;
    input \SLO_buf[25]_adj_18 ;
    output \spi_data_out_r_39__N_6114[11] ;
    input \SLO_buf[24]_adj_19 ;
    output \spi_data_out_r_39__N_6114[10] ;
    input \SLO_buf[13]_adj_20 ;
    input \SLO_buf[23]_adj_21 ;
    output \spi_data_out_r_39__N_6114[9] ;
    input \SLO_buf[4]_adj_22 ;
    input \SLO_buf[14]_adj_23 ;
    output \spi_data_out_r_39__N_5436[0] ;
    input \SLO_buf[3]_adj_24 ;
    input \SLO_buf[9]_adj_25 ;
    output \spi_data_out_r_39__N_5436[35] ;
    input \SLO_buf[2]_adj_26 ;
    input \SLO_buf[8]_adj_27 ;
    output \spi_data_out_r_39__N_6114[34] ;
    input \SLO_buf[2]_adj_28 ;
    input \SLO_buf[8]_adj_29 ;
    output \spi_data_out_r_39__N_5436[34] ;
    input \SLO_buf[1]_adj_30 ;
    input \SLO_buf[7]_adj_31 ;
    output \spi_data_out_r_39__N_5436[33] ;
    input \SLO_buf[0]_adj_32 ;
    input \SLO_buf[6]_adj_33 ;
    output \spi_data_out_r_39__N_5436[32] ;
    input \SLO_buf[12]_adj_34 ;
    input \SLO_buf[22]_adj_35 ;
    output \spi_data_out_r_39__N_6114[8] ;
    input \SLO_buf[19]_adj_36 ;
    input \SLO_buf[29]_adj_37 ;
    output \spi_data_out_r_39__N_5436[15] ;
    input \SLO_buf[18]_adj_38 ;
    input \SLO_buf[28]_adj_39 ;
    output \spi_data_out_r_39__N_5436[14] ;
    input \SLO_buf[11]_adj_40 ;
    input \SLO_buf[21]_adj_41 ;
    output \spi_data_out_r_39__N_6114[7] ;
    input \SLO_buf[10]_adj_42 ;
    input \SLO_buf[20]_adj_43 ;
    output \spi_data_out_r_39__N_6114[6] ;
    input \SLO_buf[17]_adj_44 ;
    input \SLO_buf[27]_adj_45 ;
    output \spi_data_out_r_39__N_5436[13] ;
    input \SLO_buf[16]_adj_46 ;
    input \SLO_buf[26]_adj_47 ;
    output \spi_data_out_r_39__N_5436[12] ;
    input \SLO_buf[15]_adj_48 ;
    input \SLO_buf[25]_adj_49 ;
    output \spi_data_out_r_39__N_5436[11] ;
    input \SLO_buf[1]_adj_50 ;
    input \SLO_buf[7]_adj_51 ;
    output \spi_data_out_r_39__N_6114[33] ;
    input \SLO_buf[24]_adj_52 ;
    output \spi_data_out_r_39__N_5436[10] ;
    input \SLO_buf[13]_adj_53 ;
    input \SLO_buf[23]_adj_54 ;
    output \spi_data_out_r_39__N_5436[9] ;
    output n1;
    input \SLO_buf[0]_adj_55 ;
    input \SLO_buf[6]_adj_56 ;
    output \spi_data_out_r_39__N_6114[32] ;
    input n29309;
    output n8823;
    input n29216;
    output n29205;
    input \spi_addr_r[1] ;
    input n29214;
    output n29134;
    input \SLO_buf[12]_adj_57 ;
    input \SLO_buf[22]_adj_58 ;
    output \spi_data_out_r_39__N_5436[8] ;
    input \SLO_buf[11]_adj_59 ;
    input \SLO_buf[21]_adj_60 ;
    output \spi_data_out_r_39__N_5436[7] ;
    input \SLO_buf[10]_adj_61 ;
    input \SLO_buf[20]_adj_62 ;
    output \spi_data_out_r_39__N_5436[6] ;
    output \spi_data_out_r_39__N_5436[5] ;
    output \spi_data_out_r_39__N_5436[4] ;
    output \spi_data_out_r_39__N_5436[3] ;
    output \spi_data_out_r_39__N_5436[2] ;
    input \SLO_buf[19]_adj_63 ;
    input \SLO_buf[29]_adj_64 ;
    output \spi_data_out_r_39__N_6114[15] ;
    output n1_adj_65;
    input \cs_decoded[0] ;
    output n8824;
    input \SLO_buf[5]_adj_66 ;
    output \spi_data_out_r_39__N_5436[1] ;
    output \spi_data_out_r_39__N_6114[5] ;
    output n18550;
    input \SLO_buf[18]_adj_67 ;
    output \spi_data_out_r_39__N_6114[4] ;
    input GND_net;
    input n29310;
    input \SLO_buf[4]_adj_68 ;
    input \SLO_buf[14]_adj_69 ;
    output \spi_data_out_r_39__N_5097[0] ;
    input \SLO_buf[3]_adj_70 ;
    input \SLO_buf[9]_adj_71 ;
    output \spi_data_out_r_39__N_5097[35] ;
    input \SLO_buf[2]_adj_72 ;
    input \SLO_buf[8]_adj_73 ;
    output \spi_data_out_r_39__N_5097[34] ;
    input \SLO_buf[17]_adj_74 ;
    output \spi_data_out_r_39__N_6114[3] ;
    output \spi_data_out_r_39__N_6114[2] ;
    input \SLO_buf[28]_adj_75 ;
    output \spi_data_out_r_39__N_6114[14] ;
    input mode;
    input n31;
    output n22;
    input \SLO_buf[1]_adj_76 ;
    input \SLO_buf[7]_adj_77 ;
    output \spi_data_out_r_39__N_5097[33] ;
    input \SLO_buf[0]_adj_78 ;
    input \SLO_buf[6]_adj_79 ;
    output \spi_data_out_r_39__N_5097[32] ;
    input \SLO_buf[5]_adj_80 ;
    output \spi_data_out_r_39__N_6114[1] ;
    input \SLO_buf[19]_adj_81 ;
    input \SLO_buf[29]_adj_82 ;
    output \spi_data_out_r_39__N_5097[15] ;
    input \SLO_buf[18]_adj_83 ;
    input \SLO_buf[28]_adj_84 ;
    output \spi_data_out_r_39__N_5097[14] ;
    input \SLO_buf[17]_adj_85 ;
    input \SLO_buf[27]_adj_86 ;
    output \spi_data_out_r_39__N_5097[13] ;
    input \SLO_buf[16]_adj_87 ;
    input \SLO_buf[26]_adj_88 ;
    output \spi_data_out_r_39__N_5097[12] ;
    input \SLO_buf[15]_adj_89 ;
    input \SLO_buf[25]_adj_90 ;
    output \spi_data_out_r_39__N_5097[11] ;
    input \SLO_buf[24]_adj_91 ;
    output \spi_data_out_r_39__N_5097[10] ;
    input \SLO_buf[13]_adj_92 ;
    input \SLO_buf[23]_adj_93 ;
    output \spi_data_out_r_39__N_5097[9] ;
    input \SLO_buf[12]_adj_94 ;
    input \SLO_buf[22]_adj_95 ;
    output \spi_data_out_r_39__N_5097[8] ;
    input \SLO_buf[11]_adj_96 ;
    input \SLO_buf[21]_adj_97 ;
    output \spi_data_out_r_39__N_5097[7] ;
    input \SLO_buf[10]_adj_98 ;
    input \SLO_buf[20]_adj_99 ;
    output \spi_data_out_r_39__N_5097[6] ;
    input \spi_cmd_r[1] ;
    input \spi_addr_r[0] ;
    output n29287;
    input \spi_cmd_r[0] ;
    input n29311;
    output n27286;
    input \SLO_buf[27]_adj_100 ;
    output \spi_data_out_r_39__N_6114[13] ;
    output \spi_data_out_r_39__N_5097[5] ;
    output \spi_data_out_r_39__N_5097[4] ;
    output \spi_data_out_r_39__N_5097[3] ;
    output \spi_data_out_r_39__N_5097[2] ;
    input \SLO_buf[5]_adj_101 ;
    output \spi_data_out_r_39__N_5097[1] ;
    input \SLO_buf[3]_adj_102 ;
    input \SLO_buf[9]_adj_103 ;
    output \spi_data_out_r_39__N_4419[35] ;
    input \SLO_buf[2]_adj_104 ;
    input \SLO_buf[8]_adj_105 ;
    output \spi_data_out_r_39__N_4419[34] ;
    input \SLO_buf[1]_adj_106 ;
    input \SLO_buf[7]_adj_107 ;
    output \spi_data_out_r_39__N_4419[33] ;
    input \SLO_buf[0]_adj_108 ;
    input \SLO_buf[6]_adj_109 ;
    output \spi_data_out_r_39__N_4419[32] ;
    input \SLO_buf[19]_adj_110 ;
    input \SLO_buf[29]_adj_111 ;
    output \spi_data_out_r_39__N_4419[15] ;
    input \SLO_buf[18]_adj_112 ;
    input \SLO_buf[28]_adj_113 ;
    output \spi_data_out_r_39__N_4419[14] ;
    input \SLO_buf[17]_adj_114 ;
    input \SLO_buf[27]_adj_115 ;
    output \spi_data_out_r_39__N_4419[13] ;
    input \SLO_buf[16]_adj_116 ;
    input \SLO_buf[26]_adj_117 ;
    output \spi_data_out_r_39__N_4419[12] ;
    input \SLO_buf[15]_adj_118 ;
    input \SLO_buf[25]_adj_119 ;
    output \spi_data_out_r_39__N_4419[11] ;
    input \SLO_buf[14]_adj_120 ;
    input \SLO_buf[24]_adj_121 ;
    output \spi_data_out_r_39__N_4419[10] ;
    input \SLO_buf[13]_adj_122 ;
    input \SLO_buf[23]_adj_123 ;
    output \spi_data_out_r_39__N_4419[9] ;
    input \SLO_buf[12]_adj_124 ;
    input \SLO_buf[22]_adj_125 ;
    output \spi_data_out_r_39__N_4419[8] ;
    input \SLO_buf[11]_adj_126 ;
    input \SLO_buf[21]_adj_127 ;
    output \spi_data_out_r_39__N_4419[7] ;
    input \SLO_buf[10]_adj_128 ;
    input \SLO_buf[20]_adj_129 ;
    output \spi_data_out_r_39__N_4419[6] ;
    output \spi_data_out_r_39__N_4419[5] ;
    output \spi_data_out_r_39__N_4419[4] ;
    output \spi_data_out_r_39__N_4419[3] ;
    output \spi_data_out_r_39__N_4419[2] ;
    input \SLO_buf[5]_adj_130 ;
    output \spi_data_out_r_39__N_4419[1] ;
    input \SLO_buf[4]_adj_131 ;
    output \spi_data_out_r_39__N_4419[0] ;
    input \spi_data_r[1] ;
    input \spi_data_r[2] ;
    output reset_r;
    input clk_enable_506;
    input n29106;
    output n29117;
    output n29076;
    output n29115;
    output spi_data_out_r_39__N_4490;
    output n29093;
    output n29094;
    input \spi_addr[0] ;
    input n29126;
    output clear_intrpt_N_2710;
    input \spi_cmd[1] ;
    input n29141;
    output n26933;
    input n29212;
    output n47;
    output clear_intrpt_N_2639;
    output spi_data_out_r_39__N_5507;
    output n29091;
    output n29098;
    output n29099;
    
    wire MA_Temp_N_3935 /* synthesis is_inv_clock=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    wire MA_Temp /* synthesis is_clock=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(57[5:12])
    wire clk_1MHz_derived_224 /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz_derived_224 */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire [7:0]Cnt;   // c:/s_links/sources/slot_cards/stepper.v(62[11:14])
    
    wire n29227, n28751, n29181, n11859;
    wire [51:0]SLO_buf;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    wire [51:0]SLO;   // c:/s_links/sources/slot_cards/stepper.v(63[12:15])
    
    wire clk_1MHz_derived_224_enable_46;
    wire [39:0]spi_data_out_r_39__N_4080;
    
    wire n29235, clk_1MHz_enable_98;
    wire [7:0]n199;
    wire [11:0]Cnt_NSL;   // c:/s_links/sources/slot_cards/stepper.v(61[12:19])
    wire [11:0]n1290;
    
    wire n29103, n19453, n29253, n19491, n27447, n29245, n29177, 
        spi_data_out_r_39__N_4151, n19423, clk_1MHz_enable_378, n29109, 
        n29265, n13386, NSL, clk_1MHz_derived_224_enable_27, MA_Temp_N_3949, 
        clk_1MHz_enable_99, NSL_N_4146, n29146, n24984, n29112, n24983, 
        n24982, n24981, n24980, n28750, n28752, n24979, n24978;
    wire [31:0]n153;
    
    wire n24977, n24976, n24975, n28749, MA_Temp_N_3938, n4;
    
    INV i23368 (.A(MA_Temp), .Z(MA_Temp_N_3935));
    LUT4 mux_149_i1_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[4] ), 
         .D(\SLO_buf[14] ), .Z(\spi_data_out_r_39__N_5775[0] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i1_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i36_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[3] ), 
         .D(\SLO_buf[9] ), .Z(\spi_data_out_r_39__N_5775[35] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i36_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i35_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[2] ), 
         .D(\SLO_buf[8] ), .Z(\spi_data_out_r_39__N_5775[34] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i35_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i34_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[1] ), 
         .D(\SLO_buf[7] ), .Z(\spi_data_out_r_39__N_5775[33] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i34_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i13_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29087), .C(\SLO_buf[16] ), 
         .D(\SLO_buf[26] ), .Z(\spi_data_out_r_39__N_6114[12] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i13_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i33_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[0] ), 
         .D(\SLO_buf[6] ), .Z(\spi_data_out_r_39__N_5775[32] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i33_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i16_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[19] ), 
         .D(\SLO_buf[29] ), .Z(\spi_data_out_r_39__N_5775[15] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i16_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i15_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[18] ), 
         .D(\SLO_buf[28] ), .Z(\spi_data_out_r_39__N_5775[14] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i15_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i14320_2_lut_rep_499 (.A(Cnt[4]), .B(Cnt[1]), .Z(n29227)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14320_2_lut_rep_499.init = 16'h8888;
    LUT4 n19423_bdd_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(Cnt[5]), .D(MA_Temp), 
         .Z(n28751)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;
    defparam n19423_bdd_3_lut_4_lut.init = 16'hf708;
    LUT4 mux_149_i14_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[17] ), 
         .D(\SLO_buf[27] ), .Z(\spi_data_out_r_39__N_5775[13] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i14_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(n29181), .D(Cnt[5]), 
         .Z(n11859)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff7;
    LUT4 mux_149_i13_3_lut_4_lut_adj_375 (.A(\spi_cmd[0] ), .B(n29108), 
         .C(\SLO_buf[16]_adj_11 ), .D(\SLO_buf[26]_adj_12 ), .Z(\spi_data_out_r_39__N_5775[12] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i13_3_lut_4_lut_adj_375.init = 16'hf4b0;
    LUT4 mux_149_i12_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[15] ), 
         .D(\SLO_buf[25] ), .Z(\spi_data_out_r_39__N_5775[11] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i12_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i11_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[14] ), 
         .D(\SLO_buf[24] ), .Z(\spi_data_out_r_39__N_5775[10] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i11_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i10_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[13] ), 
         .D(\SLO_buf[23] ), .Z(\spi_data_out_r_39__N_5775[9] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i10_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i9_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[12] ), 
         .D(\SLO_buf[22] ), .Z(\spi_data_out_r_39__N_5775[8] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i9_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i8_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[11] ), 
         .D(\SLO_buf[21] ), .Z(\spi_data_out_r_39__N_5775[7] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i8_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i7_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[10] ), 
         .D(\SLO_buf[20] ), .Z(\spi_data_out_r_39__N_5775[6] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i7_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i6_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[9] ), 
         .D(\SLO_buf[19] ), .Z(\spi_data_out_r_39__N_5775[5] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i6_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i5_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[8] ), 
         .D(\SLO_buf[18] ), .Z(\spi_data_out_r_39__N_5775[4] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i5_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i4_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[7] ), 
         .D(\SLO_buf[17] ), .Z(\spi_data_out_r_39__N_5775[3] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i4_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_149_i3_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[6] ), 
         .D(\SLO_buf[16]_adj_11 ), .Z(\spi_data_out_r_39__N_5775[2] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i3_3_lut_4_lut.init = 16'hf4b0;
    FD1S3AX SLO_buf_i1 (.D(SLO[0]), .CK(MA_Temp_N_3935), .Q(SLO_buf[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i1.GSR = "DISABLED";
    FD1P3AX SLO_i0 (.D(pin_io_out_8), .SP(clk_1MHz_derived_224_enable_46), 
            .CK(clk_1MHz_derived_224), .Q(SLO[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i0 (.D(spi_data_out_r_39__N_4080[0]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i0.GSR = "DISABLED";
    LUT4 mux_149_i2_3_lut_4_lut (.A(\spi_cmd[0] ), .B(n29108), .C(\SLO_buf[5] ), 
         .D(\SLO_buf[15] ), .Z(\spi_data_out_r_39__N_5775[1] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i2_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_rep_507 (.A(mode_adj_132[2]), .B(mode_adj_132[0]), .Z(n29235)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_507.init = 16'heeee;
    FD1P3IX Cnt__i0 (.D(n199[0]), .SP(clk_1MHz_enable_98), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i0.GSR = "DISABLED";
    LUT4 Select_4100_i1_2_lut_3_lut_4_lut (.A(mode_adj_132[2]), .B(mode_adj_132[0]), 
         .C(pin_io_out_9), .D(mode_adj_132[1]), .Z(\quad_b[0] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam Select_4100_i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 Select_4093_i1_2_lut_3_lut_4_lut (.A(mode_adj_132[2]), .B(mode_adj_132[0]), 
         .C(pin_io_out_8), .D(mode_adj_132[1]), .Z(\quad_a[0] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam Select_4093_i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_rep_473_3_lut (.A(mode_adj_132[2]), .B(mode_adj_132[0]), 
         .C(mode_adj_132[1]), .Z(n29201)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_473_3_lut.init = 16'hfefe;
    FD1P3IX Cnt_NSL__i0 (.D(n1290[0]), .SP(clk_1MHz_enable_55), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i0.GSR = "DISABLED";
    FD1P3IX mode__i0 (.D(n29762), .SP(clk_enable_402), .CD(n29239), .CK(clk), 
            .Q(mode_adj_132[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i0.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i11 (.D(n1290[11]), .SP(clk_1MHz_enable_55), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i11.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i10 (.D(n1290[10]), .SP(clk_1MHz_enable_55), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i10.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i9 (.D(n1290[9]), .SP(clk_1MHz_enable_55), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i9.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i8 (.D(n1290[8]), .SP(clk_1MHz_enable_55), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i8.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i7 (.D(n1290[7]), .SP(clk_1MHz_enable_55), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i7.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i6 (.D(n1290[6]), .SP(clk_1MHz_enable_55), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i6.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i5 (.D(n1290[5]), .SP(clk_1MHz_enable_55), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i5.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i4 (.D(n1290[4]), .SP(clk_1MHz_enable_55), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i4.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i3 (.D(n1290[3]), .SP(clk_1MHz_enable_55), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i3.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i2 (.D(n1290[2]), .SP(clk_1MHz_enable_55), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i2.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i1 (.D(n1290[1]), .SP(clk_1MHz_enable_55), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i1.GSR = "DISABLED";
    FD1P3IX Cnt__i7 (.D(n199[7]), .SP(clk_1MHz_enable_98), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i7.GSR = "DISABLED";
    FD1P3IX Cnt__i6 (.D(n199[6]), .SP(clk_1MHz_enable_98), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i6.GSR = "DISABLED";
    FD1P3IX Cnt__i5 (.D(n199[5]), .SP(clk_1MHz_enable_98), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i5.GSR = "DISABLED";
    FD1P3IX Cnt__i4 (.D(n199[4]), .SP(clk_1MHz_enable_98), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i4.GSR = "DISABLED";
    FD1P3IX Cnt__i3 (.D(n199[3]), .SP(clk_1MHz_enable_98), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i3.GSR = "DISABLED";
    FD1P3IX Cnt__i2 (.D(n199[2]), .SP(clk_1MHz_enable_98), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i1 (.D(n199[1]), .SP(clk_1MHz_enable_98), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i1.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i39 (.D(SLO_buf[13]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i39.GSR = "DISABLED";
    LUT4 i3_4_lut (.A(n19453), .B(Cnt[5]), .C(n29185), .D(n29253), .Z(n19491)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    FD1S3IX spi_data_out_r_i38 (.D(SLO_buf[12]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i38.GSR = "DISABLED";
    LUT4 i14513_4_lut (.A(Cnt[0]), .B(Cnt[4]), .C(n27447), .D(Cnt[1]), 
         .Z(n19453)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i14513_4_lut.init = 16'hc8c0;
    FD1S3IX spi_data_out_r_i37 (.D(SLO_buf[11]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i37.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i36 (.D(SLO_buf[10]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i36.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i35 (.D(spi_data_out_r_39__N_4080[35]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i35.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i34 (.D(spi_data_out_r_39__N_4080[34]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i34.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i33 (.D(spi_data_out_r_39__N_4080[33]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i33.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_517 (.A(\spi_addr[1] ), .B(n29761), .Z(n29245)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam i1_2_lut_rep_517.init = 16'heeee;
    LUT4 i1_2_lut_rep_449_3_lut (.A(\spi_addr[1] ), .B(n29761), .C(\spi_addr[2] ), 
         .Z(n29177)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam i1_2_lut_rep_449_3_lut.init = 16'hfefe;
    FD1S3AX spi_data_out_r_i32 (.D(spi_data_out_r_39__N_4080[32]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_376 (.A(\spi_addr[1] ), .B(n29761), .C(\spi_cmd[2] ), 
         .D(\spi_addr[2] ), .Z(n13489)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam i1_2_lut_3_lut_4_lut_adj_376.init = 16'hffef;
    LUT4 i2_3_lut_rep_450_4_lut (.A(\spi_addr[1] ), .B(n29761), .C(\spi_cmd[2] ), 
         .D(\spi_addr[2] ), .Z(n29178)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam i2_3_lut_rep_450_4_lut.init = 16'hfeff;
    FD1S3IX spi_data_out_r_i31 (.D(SLO_buf[45]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i30 (.D(SLO_buf[44]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i29 (.D(SLO_buf[43]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i28 (.D(SLO_buf[42]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i27 (.D(SLO_buf[41]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i26 (.D(SLO_buf[40]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i25 (.D(SLO_buf[39]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i24 (.D(SLO_buf[38]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i23 (.D(SLO_buf[37]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i22 (.D(SLO_buf[36]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i21 (.D(SLO_buf[35]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i20 (.D(SLO_buf[34]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i19 (.D(SLO_buf[33]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i18 (.D(SLO_buf[32]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i17 (.D(SLO_buf[31]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i16 (.D(SLO_buf[30]), .CK(clk), .CD(n29103), 
            .Q(spi_data_out_r_39__N_3818[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(spi_data_out_r_39__N_4080[15]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(spi_data_out_r_39__N_4080[14]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(spi_data_out_r_39__N_4080[13]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(spi_data_out_r_39__N_4080[12]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(spi_data_out_r_39__N_4080[11]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(spi_data_out_r_39__N_4080[10]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(spi_data_out_r_39__N_4080[9]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(spi_data_out_r_39__N_4080[8]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(spi_data_out_r_39__N_4080[7]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1P3IX digital_output_r_481 (.D(\spi_data_r[0] ), .SP(clk_enable_173), 
            .CD(n29239), .CK(clk), .Q(digital_output_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam digital_output_r_481.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_525 (.A(Cnt[7]), .B(Cnt[6]), .Z(n29253)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_rep_525.init = 16'heeee;
    LUT4 i2_3_lut_rep_453_4_lut (.A(Cnt[7]), .B(Cnt[6]), .C(Cnt[0]), .D(n27447), 
         .Z(n29181)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i2_3_lut_rep_453_4_lut.init = 16'hfffe;
    FD1S3IX i159_483 (.D(spi_data_out_r_39__N_4151), .CK(clk), .CD(n29239), 
            .Q(spi_data_out_r_39__N_3858)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam i159_483.GSR = "DISABLED";
    LUT4 mux_149_i1_3_lut_4_lut_adj_377 (.A(\spi_cmd[0] ), .B(n29087), .C(\SLO_buf[4]_adj_13 ), 
         .D(\SLO_buf[14]_adj_14 ), .Z(\spi_data_out_r_39__N_6114[0] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i1_3_lut_4_lut_adj_377.init = 16'hf4b0;
    FD1S3AX spi_data_out_r_i6 (.D(spi_data_out_r_39__N_4080[6]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(spi_data_out_r_39__N_4080[5]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(spi_data_out_r_39__N_4080[4]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(spi_data_out_r_39__N_4080[3]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(spi_data_out_r_39__N_4080[2]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(spi_data_out_r_39__N_4080[1]), .CK(clk), 
            .Q(spi_data_out_r_39__N_3818[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    LUT4 mux_149_i36_3_lut_4_lut_adj_378 (.A(\spi_cmd[0] ), .B(n29087), 
         .C(\SLO_buf[3]_adj_15 ), .D(\SLO_buf[9]_adj_16 ), .Z(\spi_data_out_r_39__N_6114[35] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i36_3_lut_4_lut_adj_378.init = 16'hf4b0;
    LUT4 i22610_2_lut_rep_409 (.A(resetn_c), .B(n19337), .Z(clk_1MHz_enable_98)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i22610_2_lut_rep_409.init = 16'hdddd;
    LUT4 i22859_2_lut_2_lut_3_lut_4_lut (.A(resetn_c), .B(n19337), .C(n19491), 
         .D(n19423), .Z(clk_1MHz_enable_378)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (C (D)))) */ ;
    defparam i22859_2_lut_2_lut_3_lut_4_lut.init = 16'h0ddd;
    LUT4 mux_149_i12_3_lut_4_lut_adj_379 (.A(\spi_cmd[0] ), .B(n29087), 
         .C(\SLO_buf[15]_adj_17 ), .D(\SLO_buf[25]_adj_18 ), .Z(\spi_data_out_r_39__N_6114[11] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i12_3_lut_4_lut_adj_379.init = 16'hf4b0;
    LUT4 mux_149_i11_3_lut_4_lut_adj_380 (.A(\spi_cmd[0] ), .B(n29087), 
         .C(\SLO_buf[14]_adj_14 ), .D(\SLO_buf[24]_adj_19 ), .Z(\spi_data_out_r_39__N_6114[10] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i11_3_lut_4_lut_adj_380.init = 16'hf4b0;
    LUT4 mux_149_i10_3_lut_4_lut_adj_381 (.A(\spi_cmd[0] ), .B(n29087), 
         .C(\SLO_buf[13]_adj_20 ), .D(\SLO_buf[23]_adj_21 ), .Z(\spi_data_out_r_39__N_6114[9] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i10_3_lut_4_lut_adj_381.init = 16'hf4b0;
    LUT4 mux_149_i1_3_lut_4_lut_adj_382 (.A(n29109), .B(n29245), .C(\SLO_buf[4]_adj_22 ), 
         .D(\SLO_buf[14]_adj_23 ), .Z(\spi_data_out_r_39__N_5436[0] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i1_3_lut_4_lut_adj_382.init = 16'hf1e0;
    LUT4 mux_149_i36_3_lut_4_lut_adj_383 (.A(n29109), .B(n29245), .C(\SLO_buf[3]_adj_24 ), 
         .D(\SLO_buf[9]_adj_25 ), .Z(\spi_data_out_r_39__N_5436[35] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i36_3_lut_4_lut_adj_383.init = 16'hf1e0;
    LUT4 mux_149_i35_3_lut_4_lut_adj_384 (.A(\spi_cmd[0] ), .B(n29087), 
         .C(\SLO_buf[2]_adj_26 ), .D(\SLO_buf[8]_adj_27 ), .Z(\spi_data_out_r_39__N_6114[34] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i35_3_lut_4_lut_adj_384.init = 16'hf4b0;
    LUT4 mux_149_i35_3_lut_4_lut_adj_385 (.A(n29109), .B(n29245), .C(\SLO_buf[2]_adj_28 ), 
         .D(\SLO_buf[8]_adj_29 ), .Z(\spi_data_out_r_39__N_5436[34] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i35_3_lut_4_lut_adj_385.init = 16'hf1e0;
    LUT4 mux_149_i34_3_lut_4_lut_adj_386 (.A(n29109), .B(n29245), .C(\SLO_buf[1]_adj_30 ), 
         .D(\SLO_buf[7]_adj_31 ), .Z(\spi_data_out_r_39__N_5436[33] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i34_3_lut_4_lut_adj_386.init = 16'hf1e0;
    LUT4 mux_149_i33_3_lut_4_lut_adj_387 (.A(n29109), .B(n29245), .C(\SLO_buf[0]_adj_32 ), 
         .D(\SLO_buf[6]_adj_33 ), .Z(\spi_data_out_r_39__N_5436[32] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i33_3_lut_4_lut_adj_387.init = 16'hf1e0;
    LUT4 mux_149_i9_3_lut_4_lut_adj_388 (.A(\spi_cmd[0] ), .B(n29087), .C(\SLO_buf[12]_adj_34 ), 
         .D(\SLO_buf[22]_adj_35 ), .Z(\spi_data_out_r_39__N_6114[8] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i9_3_lut_4_lut_adj_388.init = 16'hf4b0;
    LUT4 mux_149_i16_3_lut_4_lut_adj_389 (.A(n29109), .B(n29245), .C(\SLO_buf[19]_adj_36 ), 
         .D(\SLO_buf[29]_adj_37 ), .Z(\spi_data_out_r_39__N_5436[15] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i16_3_lut_4_lut_adj_389.init = 16'hf1e0;
    LUT4 mux_149_i15_3_lut_4_lut_adj_390 (.A(n29109), .B(n29245), .C(\SLO_buf[18]_adj_38 ), 
         .D(\SLO_buf[28]_adj_39 ), .Z(\spi_data_out_r_39__N_5436[14] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i15_3_lut_4_lut_adj_390.init = 16'hf1e0;
    LUT4 mux_149_i8_3_lut_4_lut_adj_391 (.A(\spi_cmd[0] ), .B(n29087), .C(\SLO_buf[11]_adj_40 ), 
         .D(\SLO_buf[21]_adj_41 ), .Z(\spi_data_out_r_39__N_6114[7] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i8_3_lut_4_lut_adj_391.init = 16'hf4b0;
    LUT4 mux_149_i7_3_lut_4_lut_adj_392 (.A(\spi_cmd[0] ), .B(n29087), .C(\SLO_buf[10]_adj_42 ), 
         .D(\SLO_buf[20]_adj_43 ), .Z(\spi_data_out_r_39__N_6114[6] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i7_3_lut_4_lut_adj_392.init = 16'hf4b0;
    LUT4 mux_149_i14_3_lut_4_lut_adj_393 (.A(n29109), .B(n29245), .C(\SLO_buf[17]_adj_44 ), 
         .D(\SLO_buf[27]_adj_45 ), .Z(\spi_data_out_r_39__N_5436[13] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i14_3_lut_4_lut_adj_393.init = 16'hf1e0;
    LUT4 mux_149_i13_3_lut_4_lut_adj_394 (.A(n29109), .B(n29245), .C(\SLO_buf[16]_adj_46 ), 
         .D(\SLO_buf[26]_adj_47 ), .Z(\spi_data_out_r_39__N_5436[12] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i13_3_lut_4_lut_adj_394.init = 16'hf1e0;
    LUT4 mux_149_i12_3_lut_4_lut_adj_395 (.A(n29109), .B(n29245), .C(\SLO_buf[15]_adj_48 ), 
         .D(\SLO_buf[25]_adj_49 ), .Z(\spi_data_out_r_39__N_5436[11] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i12_3_lut_4_lut_adj_395.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_537 (.A(mode_adj_132[1]), .B(mode_adj_132[2]), .Z(n29265)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(71[15:39])
    defparam i1_2_lut_rep_537.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_457_3_lut (.A(mode_adj_132[1]), .B(mode_adj_132[2]), 
         .C(mode_adj_132[0]), .Z(n29185)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(71[15:39])
    defparam i1_2_lut_rep_457_3_lut.init = 16'hbfbf;
    LUT4 mux_149_i34_3_lut_4_lut_adj_396 (.A(\spi_cmd[0] ), .B(n29087), 
         .C(\SLO_buf[1]_adj_50 ), .D(\SLO_buf[7]_adj_51 ), .Z(\spi_data_out_r_39__N_6114[33] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i34_3_lut_4_lut_adj_396.init = 16'hf4b0;
    LUT4 i1_2_lut_3_lut (.A(mode_adj_132[1]), .B(mode_adj_132[2]), .C(mode_adj_132[0]), 
         .Z(n13386)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(71[15:39])
    defparam i1_2_lut_3_lut.init = 16'hfbfb;
    LUT4 mux_149_i11_3_lut_4_lut_adj_397 (.A(n29109), .B(n29245), .C(\SLO_buf[14]_adj_23 ), 
         .D(\SLO_buf[24]_adj_52 ), .Z(\spi_data_out_r_39__N_5436[10] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i11_3_lut_4_lut_adj_397.init = 16'hf1e0;
    LUT4 mux_149_i10_3_lut_4_lut_adj_398 (.A(n29109), .B(n29245), .C(\SLO_buf[13]_adj_53 ), 
         .D(\SLO_buf[23]_adj_54 ), .Z(\spi_data_out_r_39__N_5436[9] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i10_3_lut_4_lut_adj_398.init = 16'hf1e0;
    LUT4 Select_4022_i1_2_lut_3_lut_4_lut (.A(mode_adj_132[1]), .B(mode_adj_132[2]), 
         .C(NSL), .D(mode_adj_132[0]), .Z(n1)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(71[15:39])
    defparam Select_4022_i1_2_lut_3_lut_4_lut.init = 16'h4000;
    FD1P3IX SLO_i45 (.D(SLO[44]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i45.GSR = "DISABLED";
    FD1P3IX SLO_i44 (.D(SLO[43]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i44.GSR = "DISABLED";
    FD1P3IX SLO_i43 (.D(SLO[42]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i43.GSR = "DISABLED";
    FD1P3IX SLO_i42 (.D(SLO[41]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i42.GSR = "DISABLED";
    FD1P3IX SLO_i41 (.D(SLO[40]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i41.GSR = "DISABLED";
    FD1P3IX SLO_i40 (.D(SLO[39]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i40.GSR = "DISABLED";
    FD1P3IX SLO_i39 (.D(SLO[38]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i39.GSR = "DISABLED";
    FD1P3IX SLO_i38 (.D(SLO[37]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i38.GSR = "DISABLED";
    FD1P3IX SLO_i37 (.D(SLO[36]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i37.GSR = "DISABLED";
    FD1P3IX SLO_i36 (.D(SLO[35]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i36.GSR = "DISABLED";
    FD1P3IX SLO_i35 (.D(SLO[34]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i35.GSR = "DISABLED";
    FD1P3IX SLO_i34 (.D(SLO[33]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i34.GSR = "DISABLED";
    FD1P3IX SLO_i33 (.D(SLO[32]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i33.GSR = "DISABLED";
    FD1P3IX SLO_i32 (.D(SLO[31]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i32.GSR = "DISABLED";
    FD1P3IX SLO_i31 (.D(SLO[30]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i31.GSR = "DISABLED";
    FD1P3IX SLO_i30 (.D(SLO[29]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i30.GSR = "DISABLED";
    FD1P3IX SLO_i29 (.D(SLO[28]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i29.GSR = "DISABLED";
    FD1P3IX SLO_i28 (.D(SLO[27]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i28.GSR = "DISABLED";
    FD1P3IX SLO_i27 (.D(SLO[26]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i27.GSR = "DISABLED";
    FD1P3IX SLO_i26 (.D(SLO[25]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i26.GSR = "DISABLED";
    LUT4 mux_149_i33_3_lut_4_lut_adj_399 (.A(\spi_cmd[0] ), .B(n29087), 
         .C(\SLO_buf[0]_adj_55 ), .D(\SLO_buf[6]_adj_56 ), .Z(\spi_data_out_r_39__N_6114[32] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i33_3_lut_4_lut_adj_399.init = 16'hf4b0;
    FD1P3IX SLO_i25 (.D(SLO[24]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i25.GSR = "DISABLED";
    FD1P3IX SLO_i24 (.D(SLO[23]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i24.GSR = "DISABLED";
    FD1P3IX SLO_i23 (.D(SLO[22]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i23.GSR = "DISABLED";
    FD1P3IX SLO_i22 (.D(SLO[21]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i22.GSR = "DISABLED";
    FD1P3IX SLO_i21 (.D(SLO[20]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i21.GSR = "DISABLED";
    FD1P3IX SLO_i20 (.D(SLO[19]), .SP(clk_1MHz_derived_224_enable_27), .CD(MA_Temp_N_3949), 
            .CK(clk_1MHz_derived_224), .Q(SLO[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i20.GSR = "DISABLED";
    FD1P3AX SLO_i19 (.D(SLO[18]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i19.GSR = "DISABLED";
    FD1P3AX SLO_i18 (.D(SLO[17]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i18.GSR = "DISABLED";
    FD1P3AX SLO_i17 (.D(SLO[16]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i17.GSR = "DISABLED";
    FD1P3AX SLO_i16 (.D(SLO[15]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i16.GSR = "DISABLED";
    FD1P3AX SLO_i15 (.D(SLO[14]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i15.GSR = "DISABLED";
    FD1P3AX SLO_i14 (.D(SLO[13]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i14.GSR = "DISABLED";
    FD1P3AX SLO_i13 (.D(SLO[12]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i13.GSR = "DISABLED";
    FD1P3AX SLO_i12 (.D(SLO[11]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i12.GSR = "DISABLED";
    FD1P3AX SLO_i11 (.D(SLO[10]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i11.GSR = "DISABLED";
    FD1P3AX SLO_i10 (.D(SLO[9]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i10.GSR = "DISABLED";
    FD1P3AX SLO_i9 (.D(SLO[8]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i9.GSR = "DISABLED";
    FD1P3AX SLO_i8 (.D(SLO[7]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i8.GSR = "DISABLED";
    FD1P3AX SLO_i7 (.D(SLO[6]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i7.GSR = "DISABLED";
    FD1P3AX SLO_i6 (.D(SLO[5]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i6.GSR = "DISABLED";
    FD1P3AX SLO_i5 (.D(SLO[4]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i5.GSR = "DISABLED";
    FD1P3AX SLO_i4 (.D(SLO[3]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i4.GSR = "DISABLED";
    FD1P3AX SLO_i3 (.D(SLO[2]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i3.GSR = "DISABLED";
    FD1P3AX SLO_i2 (.D(SLO[1]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i2.GSR = "DISABLED";
    FD1P3AX SLO_i1 (.D(SLO[0]), .SP(clk_1MHz_derived_224_enable_46), .CK(clk_1MHz_derived_224), 
            .Q(SLO[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i1.GSR = "DISABLED";
    FD1S3AX SLO_buf_i46 (.D(SLO[45]), .CK(MA_Temp_N_3935), .Q(SLO_buf[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i46.GSR = "DISABLED";
    FD1S3AX SLO_buf_i45 (.D(SLO[44]), .CK(MA_Temp_N_3935), .Q(SLO_buf[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i45.GSR = "DISABLED";
    FD1S3AX SLO_buf_i44 (.D(SLO[43]), .CK(MA_Temp_N_3935), .Q(SLO_buf[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i44.GSR = "DISABLED";
    FD1S3AX SLO_buf_i43 (.D(SLO[42]), .CK(MA_Temp_N_3935), .Q(SLO_buf[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i43.GSR = "DISABLED";
    FD1S3AX SLO_buf_i42 (.D(SLO[41]), .CK(MA_Temp_N_3935), .Q(SLO_buf[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i42.GSR = "DISABLED";
    FD1S3AX SLO_buf_i41 (.D(SLO[40]), .CK(MA_Temp_N_3935), .Q(SLO_buf[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i41.GSR = "DISABLED";
    FD1S3AX SLO_buf_i40 (.D(SLO[39]), .CK(MA_Temp_N_3935), .Q(SLO_buf[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i40.GSR = "DISABLED";
    FD1S3AX SLO_buf_i39 (.D(SLO[38]), .CK(MA_Temp_N_3935), .Q(SLO_buf[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i39.GSR = "DISABLED";
    FD1S3AX SLO_buf_i38 (.D(SLO[37]), .CK(MA_Temp_N_3935), .Q(SLO_buf[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i38.GSR = "DISABLED";
    FD1S3AX SLO_buf_i37 (.D(SLO[36]), .CK(MA_Temp_N_3935), .Q(SLO_buf[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i37.GSR = "DISABLED";
    FD1S3AX SLO_buf_i36 (.D(SLO[35]), .CK(MA_Temp_N_3935), .Q(SLO_buf[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i36.GSR = "DISABLED";
    FD1S3AX SLO_buf_i35 (.D(SLO[34]), .CK(MA_Temp_N_3935), .Q(SLO_buf[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i35.GSR = "DISABLED";
    FD1S3AX SLO_buf_i34 (.D(SLO[33]), .CK(MA_Temp_N_3935), .Q(SLO_buf[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i34.GSR = "DISABLED";
    FD1S3AX SLO_buf_i33 (.D(SLO[32]), .CK(MA_Temp_N_3935), .Q(SLO_buf[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i33.GSR = "DISABLED";
    FD1S3AX SLO_buf_i32 (.D(SLO[31]), .CK(MA_Temp_N_3935), .Q(SLO_buf[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i32.GSR = "DISABLED";
    FD1S3AX SLO_buf_i31 (.D(SLO[30]), .CK(MA_Temp_N_3935), .Q(SLO_buf[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i31.GSR = "DISABLED";
    FD1S3AX SLO_buf_i30 (.D(SLO[29]), .CK(MA_Temp_N_3935), .Q(SLO_buf[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i30.GSR = "DISABLED";
    LUT4 equal_91_i6_1_lut_2_lut_3_lut (.A(mode_adj_132[1]), .B(mode_adj_132[2]), 
         .C(mode_adj_132[0]), .Z(MA_Temp_N_3949)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(71[15:39])
    defparam equal_91_i6_1_lut_2_lut_3_lut.init = 16'h4040;
    LUT4 i4773_2_lut_3_lut_4_lut (.A(mode_adj_132[1]), .B(mode_adj_132[2]), 
         .C(clk_1MHz_derived_224_enable_27), .D(mode_adj_132[0]), .Z(clk_1MHz_derived_224_enable_46)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(71[15:39])
    defparam i4773_2_lut_3_lut_4_lut.init = 16'hf4f0;
    FD1S3AX SLO_buf_i29 (.D(SLO[28]), .CK(MA_Temp_N_3935), .Q(SLO_buf[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i29.GSR = "DISABLED";
    FD1S3AX SLO_buf_i28 (.D(SLO[27]), .CK(MA_Temp_N_3935), .Q(SLO_buf[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i28.GSR = "DISABLED";
    FD1S3AX SLO_buf_i27 (.D(SLO[26]), .CK(MA_Temp_N_3935), .Q(SLO_buf[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i27.GSR = "DISABLED";
    FD1S3AX SLO_buf_i26 (.D(SLO[25]), .CK(MA_Temp_N_3935), .Q(SLO_buf[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i26.GSR = "DISABLED";
    FD1S3AX SLO_buf_i25 (.D(SLO[24]), .CK(MA_Temp_N_3935), .Q(SLO_buf[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i25.GSR = "DISABLED";
    FD1S3AX SLO_buf_i24 (.D(SLO[23]), .CK(MA_Temp_N_3935), .Q(SLO_buf[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i24.GSR = "DISABLED";
    FD1S3AX SLO_buf_i23 (.D(SLO[22]), .CK(MA_Temp_N_3935), .Q(SLO_buf[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i23.GSR = "DISABLED";
    FD1S3AX SLO_buf_i22 (.D(SLO[21]), .CK(MA_Temp_N_3935), .Q(SLO_buf[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i22.GSR = "DISABLED";
    FD1S3AX SLO_buf_i21 (.D(SLO[20]), .CK(MA_Temp_N_3935), .Q(SLO_buf[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i21.GSR = "DISABLED";
    FD1S3AX SLO_buf_i20 (.D(SLO[19]), .CK(MA_Temp_N_3935), .Q(SLO_buf[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i20.GSR = "DISABLED";
    FD1S3AX SLO_buf_i19 (.D(SLO[18]), .CK(MA_Temp_N_3935), .Q(SLO_buf[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i19.GSR = "DISABLED";
    FD1S3AX SLO_buf_i18 (.D(SLO[17]), .CK(MA_Temp_N_3935), .Q(SLO_buf[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i18.GSR = "DISABLED";
    FD1S3AX SLO_buf_i17 (.D(SLO[16]), .CK(MA_Temp_N_3935), .Q(SLO_buf[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i17.GSR = "DISABLED";
    FD1S3AX SLO_buf_i16 (.D(SLO[15]), .CK(MA_Temp_N_3935), .Q(SLO_buf[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i16.GSR = "DISABLED";
    FD1S3AX SLO_buf_i15 (.D(SLO[14]), .CK(MA_Temp_N_3935), .Q(SLO_buf[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i15.GSR = "DISABLED";
    FD1S3AX SLO_buf_i14 (.D(SLO[13]), .CK(MA_Temp_N_3935), .Q(SLO_buf[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i14.GSR = "DISABLED";
    FD1S3AX SLO_buf_i13 (.D(SLO[12]), .CK(MA_Temp_N_3935), .Q(SLO_buf[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i13.GSR = "DISABLED";
    FD1S3AX SLO_buf_i12 (.D(SLO[11]), .CK(MA_Temp_N_3935), .Q(SLO_buf[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i12.GSR = "DISABLED";
    FD1S3AX SLO_buf_i11 (.D(SLO[10]), .CK(MA_Temp_N_3935), .Q(SLO_buf[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i11.GSR = "DISABLED";
    FD1S3AX SLO_buf_i10 (.D(SLO[9]), .CK(MA_Temp_N_3935), .Q(SLO_buf[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i10.GSR = "DISABLED";
    LUT4 i22699_2_lut_3_lut_3_lut_4_lut (.A(mode_adj_132[1]), .B(mode_adj_132[2]), 
         .C(mode_adj_132[0]), .D(n29309), .Z(n8823)) /* synthesis lut_function=(!(A (D)+!A (B (C+(D))+!B (D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(71[15:39])
    defparam i22699_2_lut_3_lut_3_lut_4_lut.init = 16'h00bf;
    FD1S3AX SLO_buf_i9 (.D(SLO[8]), .CK(MA_Temp_N_3935), .Q(SLO_buf[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i9.GSR = "DISABLED";
    FD1S3AX SLO_buf_i8 (.D(SLO[7]), .CK(MA_Temp_N_3935), .Q(SLO_buf[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i8.GSR = "DISABLED";
    FD1S3AX SLO_buf_i7 (.D(SLO[6]), .CK(MA_Temp_N_3935), .Q(SLO_buf[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i7.GSR = "DISABLED";
    FD1S3AX SLO_buf_i6 (.D(SLO[5]), .CK(MA_Temp_N_3935), .Q(SLO_buf[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i6.GSR = "DISABLED";
    FD1S3AX SLO_buf_i5 (.D(SLO[4]), .CK(MA_Temp_N_3935), .Q(SLO_buf[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i5.GSR = "DISABLED";
    FD1S3AX SLO_buf_i4 (.D(SLO[3]), .CK(MA_Temp_N_3935), .Q(SLO_buf[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i4.GSR = "DISABLED";
    FD1S3AX SLO_buf_i3 (.D(SLO[2]), .CK(MA_Temp_N_3935), .Q(SLO_buf[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i3.GSR = "DISABLED";
    FD1S3AX SLO_buf_i2 (.D(SLO[1]), .CK(MA_Temp_N_3935), .Q(SLO_buf[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i2.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_406_3_lut_4_lut (.A(n29216), .B(n29205), .C(\spi_addr_r[1] ), 
         .D(n29214), .Z(n29134)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_rep_406_3_lut_4_lut.init = 16'h0080;
    LUT4 mux_149_i9_3_lut_4_lut_adj_400 (.A(n29109), .B(n29245), .C(\SLO_buf[12]_adj_57 ), 
         .D(\SLO_buf[22]_adj_58 ), .Z(\spi_data_out_r_39__N_5436[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i9_3_lut_4_lut_adj_400.init = 16'hf1e0;
    LUT4 mux_149_i8_3_lut_4_lut_adj_401 (.A(n29109), .B(n29245), .C(\SLO_buf[11]_adj_59 ), 
         .D(\SLO_buf[21]_adj_60 ), .Z(\spi_data_out_r_39__N_5436[7] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i8_3_lut_4_lut_adj_401.init = 16'hf1e0;
    LUT4 mux_149_i7_3_lut_4_lut_adj_402 (.A(n29109), .B(n29245), .C(\SLO_buf[10]_adj_61 ), 
         .D(\SLO_buf[20]_adj_62 ), .Z(\spi_data_out_r_39__N_5436[6] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i7_3_lut_4_lut_adj_402.init = 16'hf1e0;
    LUT4 mux_149_i6_3_lut_4_lut_adj_403 (.A(n29109), .B(n29245), .C(\SLO_buf[9]_adj_25 ), 
         .D(\SLO_buf[19]_adj_36 ), .Z(\spi_data_out_r_39__N_5436[5] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i6_3_lut_4_lut_adj_403.init = 16'hf1e0;
    LUT4 mux_149_i5_3_lut_4_lut_adj_404 (.A(n29109), .B(n29245), .C(\SLO_buf[8]_adj_29 ), 
         .D(\SLO_buf[18]_adj_38 ), .Z(\spi_data_out_r_39__N_5436[4] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i5_3_lut_4_lut_adj_404.init = 16'hf1e0;
    LUT4 mux_149_i4_3_lut_4_lut_adj_405 (.A(n29109), .B(n29245), .C(\SLO_buf[7]_adj_31 ), 
         .D(\SLO_buf[17]_adj_44 ), .Z(\spi_data_out_r_39__N_5436[3] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i4_3_lut_4_lut_adj_405.init = 16'hf1e0;
    FD1P3AX NSL_476 (.D(NSL_N_4146), .SP(clk_1MHz_enable_99), .CK(clk_1MHz), 
            .Q(NSL)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam NSL_476.GSR = "DISABLED";
    LUT4 mux_149_i3_3_lut_4_lut_adj_406 (.A(n29109), .B(n29245), .C(\SLO_buf[6]_adj_33 ), 
         .D(\SLO_buf[16]_adj_46 ), .Z(\spi_data_out_r_39__N_5436[2] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i3_3_lut_4_lut_adj_406.init = 16'hf1e0;
    LUT4 i22622_2_lut_rep_542 (.A(MA_Temp), .B(clk_1MHz), .Z(clk_1MHz_derived_224)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[13:34])
    defparam i22622_2_lut_rep_542.init = 16'h7777;
    LUT4 i1_2_lut_rep_418_4_lut (.A(n27447), .B(Cnt[0]), .C(n29253), .D(Cnt[5]), 
         .Z(n29146)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_rep_418_4_lut.init = 16'hfffe;
    LUT4 mux_149_i16_3_lut_4_lut_adj_407 (.A(\spi_cmd[0] ), .B(n29087), 
         .C(\SLO_buf[19]_adj_63 ), .D(\SLO_buf[29]_adj_64 ), .Z(\spi_data_out_r_39__N_6114[15] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i16_3_lut_4_lut_adj_407.init = 16'hf4b0;
    LUT4 Select_4019_i1_2_lut_3_lut (.A(MA_Temp), .B(clk_1MHz), .C(mode_adj_132[2]), 
         .Z(n1_adj_65)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[13:34])
    defparam Select_4019_i1_2_lut_3_lut.init = 16'h7070;
    LUT4 Select_4042_i7_3_lut_4_lut (.A(mode_adj_132[0]), .B(n29265), .C(n29309), 
         .D(\cs_decoded[0] ), .Z(n8824)) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(71[15:39])
    defparam Select_4042_i7_3_lut_4_lut.init = 16'hf222;
    LUT4 mux_149_i2_3_lut_4_lut_adj_408 (.A(n29109), .B(n29245), .C(\SLO_buf[5]_adj_66 ), 
         .D(\SLO_buf[15]_adj_48 ), .Z(\spi_data_out_r_39__N_5436[1] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i2_3_lut_4_lut_adj_408.init = 16'hf1e0;
    LUT4 mux_149_i6_3_lut_4_lut_adj_409 (.A(\spi_cmd[0] ), .B(n29087), .C(\SLO_buf[9]_adj_16 ), 
         .D(\SLO_buf[19]_adj_63 ), .Z(\spi_data_out_r_39__N_6114[5] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i6_3_lut_4_lut_adj_409.init = 16'hf4b0;
    LUT4 i13628_2_lut (.A(\spi_cmd[2] ), .B(\spi_addr[2] ), .Z(n18550)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13628_2_lut.init = 16'h8888;
    LUT4 mux_149_i5_3_lut_4_lut_adj_410 (.A(\spi_cmd[0] ), .B(n29087), .C(\SLO_buf[8]_adj_27 ), 
         .D(\SLO_buf[18]_adj_67 ), .Z(\spi_data_out_r_39__N_6114[4] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i5_3_lut_4_lut_adj_410.init = 16'hf4b0;
    CCU2D add_551_13 (.A0(Cnt_NSL[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24984), 
          .S0(n1290[11]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_13.INIT0 = 16'h5aaa;
    defparam add_551_13.INIT1 = 16'h0000;
    defparam add_551_13.INJECT1_0 = "NO";
    defparam add_551_13.INJECT1_1 = "NO";
    LUT4 mux_149_i1_3_lut_4_lut_adj_411 (.A(n29112), .B(n29310), .C(\SLO_buf[4]_adj_68 ), 
         .D(\SLO_buf[14]_adj_69 ), .Z(\spi_data_out_r_39__N_5097[0] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i1_3_lut_4_lut_adj_411.init = 16'hf1e0;
    LUT4 mux_149_i36_3_lut_4_lut_adj_412 (.A(n29112), .B(n29310), .C(\SLO_buf[3]_adj_70 ), 
         .D(\SLO_buf[9]_adj_71 ), .Z(\spi_data_out_r_39__N_5097[35] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i36_3_lut_4_lut_adj_412.init = 16'hf1e0;
    LUT4 mux_149_i35_3_lut_4_lut_adj_413 (.A(n29112), .B(n29310), .C(\SLO_buf[2]_adj_72 ), 
         .D(\SLO_buf[8]_adj_73 ), .Z(\spi_data_out_r_39__N_5097[34] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i35_3_lut_4_lut_adj_413.init = 16'hf1e0;
    CCU2D add_551_11 (.A0(Cnt_NSL[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24983), .COUT(n24984), .S0(n1290[9]), .S1(n1290[10]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_11.INIT0 = 16'h5aaa;
    defparam add_551_11.INIT1 = 16'h5aaa;
    defparam add_551_11.INJECT1_0 = "NO";
    defparam add_551_11.INJECT1_1 = "NO";
    CCU2D add_551_9 (.A0(Cnt_NSL[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24982), .COUT(n24983), .S0(n1290[7]), .S1(n1290[8]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_9.INIT0 = 16'h5aaa;
    defparam add_551_9.INIT1 = 16'h5aaa;
    defparam add_551_9.INJECT1_0 = "NO";
    defparam add_551_9.INJECT1_1 = "NO";
    CCU2D add_551_7 (.A0(Cnt_NSL[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24981), .COUT(n24982), .S0(n1290[5]), .S1(n1290[6]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_7.INIT0 = 16'h5aaa;
    defparam add_551_7.INIT1 = 16'h5aaa;
    defparam add_551_7.INJECT1_0 = "NO";
    defparam add_551_7.INJECT1_1 = "NO";
    CCU2D add_551_5 (.A0(Cnt_NSL[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24980), .COUT(n24981), .S0(n1290[3]), .S1(n1290[4]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_5.INIT0 = 16'h5aaa;
    defparam add_551_5.INIT1 = 16'h5aaa;
    defparam add_551_5.INJECT1_0 = "NO";
    defparam add_551_5.INJECT1_1 = "NO";
    LUT4 mux_149_i4_3_lut_4_lut_adj_414 (.A(\spi_cmd[0] ), .B(n29087), .C(\SLO_buf[7]_adj_51 ), 
         .D(\SLO_buf[17]_adj_74 ), .Z(\spi_data_out_r_39__N_6114[3] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i4_3_lut_4_lut_adj_414.init = 16'hf4b0;
    LUT4 mux_149_i3_3_lut_4_lut_adj_415 (.A(\spi_cmd[0] ), .B(n29087), .C(\SLO_buf[6]_adj_56 ), 
         .D(\SLO_buf[16] ), .Z(\spi_data_out_r_39__N_6114[2] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i3_3_lut_4_lut_adj_415.init = 16'hf4b0;
    LUT4 mux_149_i15_3_lut_4_lut_adj_416 (.A(\spi_cmd[0] ), .B(n29087), 
         .C(\SLO_buf[18]_adj_67 ), .D(\SLO_buf[28]_adj_75 ), .Z(\spi_data_out_r_39__N_6114[14] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i15_3_lut_4_lut_adj_416.init = 16'hf4b0;
    LUT4 i3_3_lut_4_lut (.A(mode_adj_132[1]), .B(n29235), .C(mode), .D(n31), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_3_lut_4_lut.init = 16'hfffe;
    PFUMX i23055 (.BLUT(n28751), .ALUT(n28750), .C0(n19491), .Z(n28752));
    CCU2D add_551_3 (.A0(Cnt_NSL[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24979), .COUT(n24980), .S0(n1290[1]), .S1(n1290[2]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_3.INIT0 = 16'h5aaa;
    defparam add_551_3.INIT1 = 16'h5aaa;
    defparam add_551_3.INJECT1_0 = "NO";
    defparam add_551_3.INJECT1_1 = "NO";
    CCU2D add_551_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24979), .S1(n1290[0]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_1.INIT0 = 16'hF000;
    defparam add_551_1.INIT1 = 16'h5555;
    defparam add_551_1.INJECT1_0 = "NO";
    defparam add_551_1.INJECT1_1 = "NO";
    CCU2D add_552_9 (.A0(Cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24978), 
          .S0(n153[7]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_9.INIT0 = 16'h5aaa;
    defparam add_552_9.INIT1 = 16'h0000;
    defparam add_552_9.INJECT1_0 = "NO";
    defparam add_552_9.INJECT1_1 = "NO";
    CCU2D add_552_7 (.A0(Cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24977), 
          .COUT(n24978), .S0(n153[5]), .S1(n153[6]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_7.INIT0 = 16'h5aaa;
    defparam add_552_7.INIT1 = 16'h5aaa;
    defparam add_552_7.INJECT1_0 = "NO";
    defparam add_552_7.INJECT1_1 = "NO";
    LUT4 mux_149_i34_3_lut_4_lut_adj_417 (.A(n29112), .B(n29310), .C(\SLO_buf[1]_adj_76 ), 
         .D(\SLO_buf[7]_adj_77 ), .Z(\spi_data_out_r_39__N_5097[33] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i34_3_lut_4_lut_adj_417.init = 16'hf1e0;
    LUT4 mux_149_i33_3_lut_4_lut_adj_418 (.A(n29112), .B(n29310), .C(\SLO_buf[0]_adj_78 ), 
         .D(\SLO_buf[6]_adj_79 ), .Z(\spi_data_out_r_39__N_5097[32] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i33_3_lut_4_lut_adj_418.init = 16'hf1e0;
    CCU2D add_552_5 (.A0(Cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24976), 
          .COUT(n24977), .S0(n153[3]), .S1(n153[4]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_5.INIT0 = 16'h5aaa;
    defparam add_552_5.INIT1 = 16'h5aaa;
    defparam add_552_5.INJECT1_0 = "NO";
    defparam add_552_5.INJECT1_1 = "NO";
    CCU2D add_552_3 (.A0(Cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24975), 
          .COUT(n24976), .S0(n153[1]), .S1(n153[2]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_3.INIT0 = 16'h5aaa;
    defparam add_552_3.INIT1 = 16'h5aaa;
    defparam add_552_3.INJECT1_0 = "NO";
    defparam add_552_3.INJECT1_1 = "NO";
    CCU2D add_552_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24975), 
          .S1(n153[0]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_1.INIT0 = 16'hF000;
    defparam add_552_1.INIT1 = 16'h5555;
    defparam add_552_1.INJECT1_0 = "NO";
    defparam add_552_1.INJECT1_1 = "NO";
    LUT4 mux_149_i2_3_lut_4_lut_adj_419 (.A(\spi_cmd[0] ), .B(n29087), .C(\SLO_buf[5]_adj_80 ), 
         .D(\SLO_buf[15]_adj_17 ), .Z(\spi_data_out_r_39__N_6114[1] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i2_3_lut_4_lut_adj_419.init = 16'hf4b0;
    LUT4 mux_149_i16_3_lut_4_lut_adj_420 (.A(n29112), .B(n29310), .C(\SLO_buf[19]_adj_81 ), 
         .D(\SLO_buf[29]_adj_82 ), .Z(\spi_data_out_r_39__N_5097[15] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i16_3_lut_4_lut_adj_420.init = 16'hf1e0;
    LUT4 mux_149_i15_3_lut_4_lut_adj_421 (.A(n29112), .B(n29310), .C(\SLO_buf[18]_adj_83 ), 
         .D(\SLO_buf[28]_adj_84 ), .Z(\spi_data_out_r_39__N_5097[14] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i15_3_lut_4_lut_adj_421.init = 16'hf1e0;
    LUT4 mux_149_i14_3_lut_4_lut_adj_422 (.A(n29112), .B(n29310), .C(\SLO_buf[17]_adj_85 ), 
         .D(\SLO_buf[27]_adj_86 ), .Z(\spi_data_out_r_39__N_5097[13] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i14_3_lut_4_lut_adj_422.init = 16'hf1e0;
    LUT4 mux_149_i13_3_lut_4_lut_adj_423 (.A(n29112), .B(n29310), .C(\SLO_buf[16]_adj_87 ), 
         .D(\SLO_buf[26]_adj_88 ), .Z(\spi_data_out_r_39__N_5097[12] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i13_3_lut_4_lut_adj_423.init = 16'hf1e0;
    LUT4 mux_149_i12_3_lut_4_lut_adj_424 (.A(n29112), .B(n29310), .C(\SLO_buf[15]_adj_89 ), 
         .D(\SLO_buf[25]_adj_90 ), .Z(\spi_data_out_r_39__N_5097[11] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i12_3_lut_4_lut_adj_424.init = 16'hf1e0;
    LUT4 mux_149_i11_3_lut_4_lut_adj_425 (.A(n29112), .B(n29310), .C(\SLO_buf[14]_adj_69 ), 
         .D(\SLO_buf[24]_adj_91 ), .Z(\spi_data_out_r_39__N_5097[10] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i11_3_lut_4_lut_adj_425.init = 16'hf1e0;
    LUT4 mux_149_i10_3_lut_4_lut_adj_426 (.A(n29112), .B(n29310), .C(\SLO_buf[13]_adj_92 ), 
         .D(\SLO_buf[23]_adj_93 ), .Z(\spi_data_out_r_39__N_5097[9] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i10_3_lut_4_lut_adj_426.init = 16'hf1e0;
    LUT4 mux_149_i9_3_lut_4_lut_adj_427 (.A(n29112), .B(n29310), .C(\SLO_buf[12]_adj_94 ), 
         .D(\SLO_buf[22]_adj_95 ), .Z(\spi_data_out_r_39__N_5097[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i9_3_lut_4_lut_adj_427.init = 16'hf1e0;
    LUT4 mux_149_i8_3_lut_4_lut_adj_428 (.A(n29112), .B(n29310), .C(\SLO_buf[11]_adj_96 ), 
         .D(\SLO_buf[21]_adj_97 ), .Z(\spi_data_out_r_39__N_5097[7] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i8_3_lut_4_lut_adj_428.init = 16'hf1e0;
    LUT4 mux_149_i7_3_lut_4_lut_adj_429 (.A(n29112), .B(n29310), .C(\SLO_buf[10]_adj_98 ), 
         .D(\SLO_buf[20]_adj_99 ), .Z(\spi_data_out_r_39__N_5097[6] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i7_3_lut_4_lut_adj_429.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_559 (.A(\spi_cmd_r[1] ), .B(\spi_addr_r[0] ), .Z(n29287)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_559.init = 16'h2222;
    LUT4 i1_2_lut_rep_477_3_lut (.A(\spi_cmd_r[1] ), .B(\spi_addr_r[0] ), 
         .C(\spi_cmd_r[0] ), .Z(n29205)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam i1_2_lut_rep_477_3_lut.init = 16'h0202;
    LUT4 i1_2_lut_3_lut_4_lut_adj_430 (.A(\spi_cmd_r[1] ), .B(\spi_addr_r[0] ), 
         .C(n29311), .D(\spi_cmd_r[0] ), .Z(n27286)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_430.init = 16'h2000;
    LUT4 mux_149_i14_3_lut_4_lut_adj_431 (.A(\spi_cmd[0] ), .B(n29087), 
         .C(\SLO_buf[17]_adj_74 ), .D(\SLO_buf[27]_adj_100 ), .Z(\spi_data_out_r_39__N_6114[13] )) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i14_3_lut_4_lut_adj_431.init = 16'hf4b0;
    LUT4 mux_149_i6_3_lut_4_lut_adj_432 (.A(n29112), .B(n29310), .C(\SLO_buf[9]_adj_71 ), 
         .D(\SLO_buf[19]_adj_81 ), .Z(\spi_data_out_r_39__N_5097[5] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i6_3_lut_4_lut_adj_432.init = 16'hf1e0;
    LUT4 mux_149_i5_3_lut_4_lut_adj_433 (.A(n29112), .B(n29310), .C(\SLO_buf[8]_adj_73 ), 
         .D(\SLO_buf[18]_adj_83 ), .Z(\spi_data_out_r_39__N_5097[4] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i5_3_lut_4_lut_adj_433.init = 16'hf1e0;
    LUT4 mux_149_i4_3_lut_4_lut_adj_434 (.A(n29112), .B(n29310), .C(\SLO_buf[7]_adj_77 ), 
         .D(\SLO_buf[17]_adj_85 ), .Z(\spi_data_out_r_39__N_5097[3] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i4_3_lut_4_lut_adj_434.init = 16'hf1e0;
    LUT4 mux_149_i3_3_lut_4_lut_adj_435 (.A(n29112), .B(n29310), .C(\SLO_buf[6]_adj_79 ), 
         .D(\SLO_buf[16]_adj_87 ), .Z(\spi_data_out_r_39__N_5097[2] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i3_3_lut_4_lut_adj_435.init = 16'hf1e0;
    LUT4 mux_149_i2_3_lut_4_lut_adj_436 (.A(n29112), .B(n29310), .C(\SLO_buf[5]_adj_101 ), 
         .D(\SLO_buf[15]_adj_89 ), .Z(\spi_data_out_r_39__N_5097[1] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i2_3_lut_4_lut_adj_436.init = 16'hf1e0;
    LUT4 mux_149_i36_3_lut_4_lut_adj_437 (.A(n29112), .B(n29245), .C(\SLO_buf[3]_adj_102 ), 
         .D(\SLO_buf[9]_adj_103 ), .Z(\spi_data_out_r_39__N_4419[35] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i36_3_lut_4_lut_adj_437.init = 16'hf1e0;
    LUT4 mux_149_i35_3_lut_4_lut_adj_438 (.A(n29112), .B(n29245), .C(\SLO_buf[2]_adj_104 ), 
         .D(\SLO_buf[8]_adj_105 ), .Z(\spi_data_out_r_39__N_4419[34] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i35_3_lut_4_lut_adj_438.init = 16'hf1e0;
    LUT4 mux_149_i34_3_lut_4_lut_adj_439 (.A(n29112), .B(n29245), .C(\SLO_buf[1]_adj_106 ), 
         .D(\SLO_buf[7]_adj_107 ), .Z(\spi_data_out_r_39__N_4419[33] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i34_3_lut_4_lut_adj_439.init = 16'hf1e0;
    LUT4 mux_149_i33_3_lut_4_lut_adj_440 (.A(n29112), .B(n29245), .C(\SLO_buf[0]_adj_108 ), 
         .D(\SLO_buf[6]_adj_109 ), .Z(\spi_data_out_r_39__N_4419[32] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i33_3_lut_4_lut_adj_440.init = 16'hf1e0;
    LUT4 mux_149_i16_3_lut_4_lut_adj_441 (.A(n29112), .B(n29245), .C(\SLO_buf[19]_adj_110 ), 
         .D(\SLO_buf[29]_adj_111 ), .Z(\spi_data_out_r_39__N_4419[15] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i16_3_lut_4_lut_adj_441.init = 16'hf1e0;
    LUT4 mux_149_i15_3_lut_4_lut_adj_442 (.A(n29112), .B(n29245), .C(\SLO_buf[18]_adj_112 ), 
         .D(\SLO_buf[28]_adj_113 ), .Z(\spi_data_out_r_39__N_4419[14] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i15_3_lut_4_lut_adj_442.init = 16'hf1e0;
    LUT4 mux_149_i14_3_lut_4_lut_adj_443 (.A(n29112), .B(n29245), .C(\SLO_buf[17]_adj_114 ), 
         .D(\SLO_buf[27]_adj_115 ), .Z(\spi_data_out_r_39__N_4419[13] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i14_3_lut_4_lut_adj_443.init = 16'hf1e0;
    LUT4 mux_149_i13_3_lut_4_lut_adj_444 (.A(n29112), .B(n29245), .C(\SLO_buf[16]_adj_116 ), 
         .D(\SLO_buf[26]_adj_117 ), .Z(\spi_data_out_r_39__N_4419[12] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i13_3_lut_4_lut_adj_444.init = 16'hf1e0;
    LUT4 mux_149_i12_3_lut_4_lut_adj_445 (.A(n29112), .B(n29245), .C(\SLO_buf[15]_adj_118 ), 
         .D(\SLO_buf[25]_adj_119 ), .Z(\spi_data_out_r_39__N_4419[11] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i12_3_lut_4_lut_adj_445.init = 16'hf1e0;
    LUT4 mux_149_i11_3_lut_4_lut_adj_446 (.A(n29112), .B(n29245), .C(\SLO_buf[14]_adj_120 ), 
         .D(\SLO_buf[24]_adj_121 ), .Z(\spi_data_out_r_39__N_4419[10] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i11_3_lut_4_lut_adj_446.init = 16'hf1e0;
    LUT4 mux_149_i10_3_lut_4_lut_adj_447 (.A(n29112), .B(n29245), .C(\SLO_buf[13]_adj_122 ), 
         .D(\SLO_buf[23]_adj_123 ), .Z(\spi_data_out_r_39__N_4419[9] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i10_3_lut_4_lut_adj_447.init = 16'hf1e0;
    LUT4 mux_149_i9_3_lut_4_lut_adj_448 (.A(n29112), .B(n29245), .C(\SLO_buf[12]_adj_124 ), 
         .D(\SLO_buf[22]_adj_125 ), .Z(\spi_data_out_r_39__N_4419[8] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i9_3_lut_4_lut_adj_448.init = 16'hf1e0;
    LUT4 mux_149_i8_3_lut_4_lut_adj_449 (.A(n29112), .B(n29245), .C(\SLO_buf[11]_adj_126 ), 
         .D(\SLO_buf[21]_adj_127 ), .Z(\spi_data_out_r_39__N_4419[7] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i8_3_lut_4_lut_adj_449.init = 16'hf1e0;
    LUT4 mux_149_i7_3_lut_4_lut_adj_450 (.A(n29112), .B(n29245), .C(\SLO_buf[10]_adj_128 ), 
         .D(\SLO_buf[20]_adj_129 ), .Z(\spi_data_out_r_39__N_4419[6] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i7_3_lut_4_lut_adj_450.init = 16'hf1e0;
    LUT4 mux_149_i6_3_lut_4_lut_adj_451 (.A(n29112), .B(n29245), .C(\SLO_buf[9]_adj_103 ), 
         .D(\SLO_buf[19]_adj_110 ), .Z(\spi_data_out_r_39__N_4419[5] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i6_3_lut_4_lut_adj_451.init = 16'hf1e0;
    LUT4 mux_149_i5_3_lut_4_lut_adj_452 (.A(n29112), .B(n29245), .C(\SLO_buf[8]_adj_105 ), 
         .D(\SLO_buf[18]_adj_112 ), .Z(\spi_data_out_r_39__N_4419[4] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i5_3_lut_4_lut_adj_452.init = 16'hf1e0;
    LUT4 mux_149_i4_3_lut_4_lut_adj_453 (.A(n29112), .B(n29245), .C(\SLO_buf[7]_adj_107 ), 
         .D(\SLO_buf[17]_adj_114 ), .Z(\spi_data_out_r_39__N_4419[3] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i4_3_lut_4_lut_adj_453.init = 16'hf1e0;
    LUT4 mux_149_i3_3_lut_4_lut_adj_454 (.A(n29112), .B(n29245), .C(\SLO_buf[6]_adj_109 ), 
         .D(\SLO_buf[16]_adj_116 ), .Z(\spi_data_out_r_39__N_4419[2] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i3_3_lut_4_lut_adj_454.init = 16'hf1e0;
    LUT4 mux_149_i2_3_lut_4_lut_adj_455 (.A(n29112), .B(n29245), .C(\SLO_buf[5]_adj_130 ), 
         .D(\SLO_buf[15]_adj_118 ), .Z(\spi_data_out_r_39__N_4419[1] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i2_3_lut_4_lut_adj_455.init = 16'hf1e0;
    LUT4 mux_149_i1_3_lut_4_lut_adj_456 (.A(n29112), .B(n29245), .C(\SLO_buf[4]_adj_131 ), 
         .D(\SLO_buf[14]_adj_120 ), .Z(\spi_data_out_r_39__N_4419[0] )) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i1_3_lut_4_lut_adj_456.init = 16'hf1e0;
    LUT4 i117_4_lut (.A(n29146), .B(n13386), .C(Cnt[4]), .D(Cnt[1]), 
         .Z(clk_1MHz_derived_224_enable_27)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(132[15:49])
    defparam i117_4_lut.init = 16'h3332;
    FD1P3IX mode__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_402), .CD(n29239), 
            .CK(clk), .Q(mode_adj_132[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i1.GSR = "DISABLED";
    FD1P3IX mode__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_402), .CD(n29239), 
            .CK(clk), .Q(mode_adj_132[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i2.GSR = "DISABLED";
    FD1P3IX reset_r_480 (.D(n29106), .SP(clk_enable_506), .CD(n29239), 
            .CK(clk), .Q(reset_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam reset_r_480.GSR = "DISABLED";
    LUT4 mux_149_i1_3_lut_4_lut_adj_457 (.A(n13489), .B(n29117), .C(SLO_buf[4]), 
         .D(SLO_buf[14]), .Z(spi_data_out_r_39__N_4080[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i1_3_lut_4_lut_adj_457.init = 16'hf1e0;
    LUT4 mux_149_i36_3_lut_4_lut_adj_458 (.A(n13489), .B(n29117), .C(SLO_buf[3]), 
         .D(SLO_buf[9]), .Z(spi_data_out_r_39__N_4080[35])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i36_3_lut_4_lut_adj_458.init = 16'hf1e0;
    LUT4 mux_149_i35_3_lut_4_lut_adj_459 (.A(n13489), .B(n29117), .C(SLO_buf[2]), 
         .D(SLO_buf[8]), .Z(spi_data_out_r_39__N_4080[34])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i35_3_lut_4_lut_adj_459.init = 16'hf1e0;
    LUT4 mux_149_i34_3_lut_4_lut_adj_460 (.A(n13489), .B(n29117), .C(SLO_buf[1]), 
         .D(SLO_buf[7]), .Z(spi_data_out_r_39__N_4080[33])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i34_3_lut_4_lut_adj_460.init = 16'hf1e0;
    LUT4 mux_149_i33_3_lut_4_lut_adj_461 (.A(n13489), .B(n29117), .C(SLO_buf[0]), 
         .D(SLO_buf[6]), .Z(spi_data_out_r_39__N_4080[32])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i33_3_lut_4_lut_adj_461.init = 16'hf1e0;
    LUT4 mux_149_i16_3_lut_4_lut_adj_462 (.A(n13489), .B(n29117), .C(SLO_buf[19]), 
         .D(SLO_buf[29]), .Z(spi_data_out_r_39__N_4080[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i16_3_lut_4_lut_adj_462.init = 16'hf1e0;
    LUT4 mux_149_i15_3_lut_4_lut_adj_463 (.A(n13489), .B(n29117), .C(SLO_buf[18]), 
         .D(SLO_buf[28]), .Z(spi_data_out_r_39__N_4080[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i15_3_lut_4_lut_adj_463.init = 16'hf1e0;
    LUT4 mux_149_i14_3_lut_4_lut_adj_464 (.A(n13489), .B(n29117), .C(SLO_buf[17]), 
         .D(SLO_buf[27]), .Z(spi_data_out_r_39__N_4080[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i14_3_lut_4_lut_adj_464.init = 16'hf1e0;
    LUT4 mux_149_i13_3_lut_4_lut_adj_465 (.A(n13489), .B(n29117), .C(SLO_buf[16]), 
         .D(SLO_buf[26]), .Z(spi_data_out_r_39__N_4080[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i13_3_lut_4_lut_adj_465.init = 16'hf1e0;
    LUT4 mux_149_i12_3_lut_4_lut_adj_466 (.A(n13489), .B(n29117), .C(SLO_buf[15]), 
         .D(SLO_buf[25]), .Z(spi_data_out_r_39__N_4080[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i12_3_lut_4_lut_adj_466.init = 16'hf1e0;
    LUT4 mux_149_i11_3_lut_4_lut_adj_467 (.A(n13489), .B(n29117), .C(SLO_buf[14]), 
         .D(SLO_buf[24]), .Z(spi_data_out_r_39__N_4080[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i11_3_lut_4_lut_adj_467.init = 16'hf1e0;
    LUT4 mux_149_i10_3_lut_4_lut_adj_468 (.A(n13489), .B(n29117), .C(SLO_buf[13]), 
         .D(SLO_buf[23]), .Z(spi_data_out_r_39__N_4080[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i10_3_lut_4_lut_adj_468.init = 16'hf1e0;
    LUT4 mux_149_i9_3_lut_4_lut_adj_469 (.A(n13489), .B(n29117), .C(SLO_buf[12]), 
         .D(SLO_buf[22]), .Z(spi_data_out_r_39__N_4080[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i9_3_lut_4_lut_adj_469.init = 16'hf1e0;
    LUT4 mux_149_i8_3_lut_4_lut_adj_470 (.A(n13489), .B(n29117), .C(SLO_buf[11]), 
         .D(SLO_buf[21]), .Z(spi_data_out_r_39__N_4080[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i8_3_lut_4_lut_adj_470.init = 16'hf1e0;
    LUT4 mux_149_i7_3_lut_4_lut_adj_471 (.A(n13489), .B(n29117), .C(SLO_buf[10]), 
         .D(SLO_buf[20]), .Z(spi_data_out_r_39__N_4080[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i7_3_lut_4_lut_adj_471.init = 16'hf1e0;
    LUT4 mux_149_i6_3_lut_4_lut_adj_472 (.A(n13489), .B(n29117), .C(SLO_buf[9]), 
         .D(SLO_buf[19]), .Z(spi_data_out_r_39__N_4080[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i6_3_lut_4_lut_adj_472.init = 16'hf1e0;
    LUT4 mux_149_i5_3_lut_4_lut_adj_473 (.A(n13489), .B(n29117), .C(SLO_buf[8]), 
         .D(SLO_buf[18]), .Z(spi_data_out_r_39__N_4080[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i5_3_lut_4_lut_adj_473.init = 16'hf1e0;
    LUT4 mux_149_i4_3_lut_4_lut_adj_474 (.A(n13489), .B(n29117), .C(SLO_buf[7]), 
         .D(SLO_buf[17]), .Z(spi_data_out_r_39__N_4080[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i4_3_lut_4_lut_adj_474.init = 16'hf1e0;
    LUT4 mux_149_i3_3_lut_4_lut_adj_475 (.A(n13489), .B(n29117), .C(SLO_buf[6]), 
         .D(SLO_buf[16]), .Z(spi_data_out_r_39__N_4080[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i3_3_lut_4_lut_adj_475.init = 16'hf1e0;
    LUT4 mux_149_i2_3_lut_4_lut_adj_476 (.A(n13489), .B(n29117), .C(SLO_buf[5]), 
         .D(SLO_buf[15]), .Z(spi_data_out_r_39__N_4080[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam mux_149_i2_3_lut_4_lut_adj_476.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_348_3_lut_4_lut (.A(n29117), .B(n18550), .C(\spi_cmd[0] ), 
         .D(\spi_addr[1] ), .Z(n29076)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(202[15:42])
    defparam i1_2_lut_rep_348_3_lut_4_lut.init = 16'hfbff;
    LUT4 i22632_2_lut_4_lut (.A(\spi_addr[2] ), .B(n29115), .C(\spi_cmd[2] ), 
         .D(\spi_addr[1] ), .Z(spi_data_out_r_39__N_4490)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i22632_2_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_365_4_lut (.A(\spi_addr[2] ), .B(n29115), .C(\spi_cmd[2] ), 
         .D(n29310), .Z(n29093)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i1_2_lut_rep_365_4_lut.init = 16'hffef;
    LUT4 i1_2_lut_rep_366_4_lut (.A(\spi_addr[2] ), .B(n29115), .C(\spi_cmd[2] ), 
         .D(n29245), .Z(n29094)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i1_2_lut_rep_366_4_lut.init = 16'hffef;
    LUT4 n28752_bdd_3_lut (.A(n28752), .B(n28749), .C(n29181), .Z(MA_Temp_N_3938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28752_bdd_3_lut.init = 16'hcaca;
    LUT4 i22924_2_lut_2_lut_3_lut_4_lut (.A(\spi_addr[0] ), .B(n29126), 
         .C(n29177), .D(\spi_cmd[2] ), .Z(clear_intrpt_N_2710)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i22924_2_lut_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i22669_3_lut_rep_380_4_lut (.A(\spi_addr[0] ), .B(n29126), .C(\spi_addr[1] ), 
         .D(n18550), .Z(n29108)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i22669_3_lut_rep_380_4_lut.init = 16'h0200;
    LUT4 i2_3_lut_rep_384_4_lut (.A(\spi_addr[0] ), .B(n29126), .C(\spi_cmd[2] ), 
         .D(\spi_addr[2] ), .Z(n29112)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i2_3_lut_rep_384_4_lut.init = 16'hffdf;
    LUT4 n19423_bdd_4_lut_23250 (.A(n19423), .B(n29227), .C(MA_Temp), 
         .D(Cnt[5]), .Z(n28750)) /* synthesis lut_function=(!(A+(B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam n19423_bdd_4_lut_23250.init = 16'h1450;
    LUT4 n19423_bdd_3_lut_23054 (.A(n19423), .B(n19491), .C(MA_Temp), 
         .Z(n28749)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam n19423_bdd_3_lut_23054.init = 16'h7070;
    LUT4 i1_2_lut (.A(Cnt[2]), .B(Cnt[3]), .Z(n27447)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i2_3_lut (.A(\spi_cmd[1] ), .B(n29141), .C(\spi_cmd[2] ), .Z(n26933)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i2_3_lut.init = 16'hefef;
    LUT4 i2_3_lut_4_lut (.A(\spi_addr[0] ), .B(n29126), .C(\spi_cmd[2] ), 
         .D(n29212), .Z(n47)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i2_3_lut_4_lut.init = 16'hffef;
    LUT4 i22927_2_lut_2_lut_3_lut_4_lut (.A(\spi_addr[0] ), .B(n29126), 
         .C(n29177), .D(\spi_cmd[2] ), .Z(clear_intrpt_N_2639)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i22927_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 i22678_2_lut_rep_359_3_lut_4_lut (.A(\spi_addr[0] ), .B(n29126), 
         .C(\spi_addr[1] ), .D(n18550), .Z(n29087)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i22678_2_lut_rep_359_3_lut_4_lut.init = 16'h1000;
    LUT4 i22659_2_lut_3_lut_4_lut (.A(\spi_addr[0] ), .B(n29126), .C(\spi_addr[1] ), 
         .D(n18550), .Z(spi_data_out_r_39__N_5507)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i22659_2_lut_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_2_lut_rep_363_3_lut_4_lut (.A(\spi_addr[0] ), .B(n29126), .C(n29245), 
         .D(n18550), .Z(n29091)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i1_2_lut_rep_363_3_lut_4_lut.init = 16'hfeff;
    LUT4 i2_4_lut (.A(n29117), .B(\spi_addr[1] ), .C(\spi_cmd[2] ), .D(\spi_addr[2] ), 
         .Z(spi_data_out_r_39__N_4151)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_4_lut.init = 16'h0010;
    LUT4 i2_4_lut_adj_477 (.A(Cnt_NSL[11]), .B(Cnt_NSL[9]), .C(Cnt_NSL[10]), 
         .D(n4), .Z(n19337)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_477.init = 16'ha080;
    LUT4 i13630_2_lut_3_lut (.A(n19423), .B(n19491), .C(n153[0]), .Z(n199[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13630_2_lut_3_lut.init = 16'h7070;
    LUT4 i13835_2_lut_3_lut (.A(n19423), .B(n19491), .C(n153[7]), .Z(n199[7])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13835_2_lut_3_lut.init = 16'h7070;
    LUT4 i13836_2_lut_3_lut (.A(n19423), .B(n19491), .C(n153[6]), .Z(n199[6])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13836_2_lut_3_lut.init = 16'h7070;
    LUT4 i13837_2_lut_3_lut (.A(n19423), .B(n19491), .C(n153[5]), .Z(n199[5])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13837_2_lut_3_lut.init = 16'h7070;
    LUT4 i13838_2_lut_3_lut (.A(n19423), .B(n19491), .C(n153[4]), .Z(n199[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13838_2_lut_3_lut.init = 16'h7070;
    LUT4 i13839_2_lut_3_lut (.A(n19423), .B(n19491), .C(n153[3]), .Z(n199[3])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13839_2_lut_3_lut.init = 16'h7070;
    LUT4 i13840_2_lut_3_lut (.A(n19423), .B(n19491), .C(n153[2]), .Z(n199[2])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13840_2_lut_3_lut.init = 16'h7070;
    LUT4 i13841_2_lut_3_lut (.A(n19423), .B(n19491), .C(n153[1]), .Z(n199[1])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13841_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_387_3_lut (.A(\spi_cmd[1] ), .B(n29141), .C(\spi_addr[0] ), 
         .Z(n29115)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i1_2_lut_rep_387_3_lut.init = 16'hdfdf;
    LUT4 i1_2_lut_rep_370_3_lut_4_lut (.A(\spi_cmd[1] ), .B(n29141), .C(\spi_cmd[2] ), 
         .D(\spi_addr[0] ), .Z(n29098)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i1_2_lut_rep_370_3_lut_4_lut.init = 16'hfdff;
    LUT4 i1_2_lut_rep_389_3_lut (.A(\spi_cmd[1] ), .B(n29141), .C(\spi_addr[0] ), 
         .Z(n29117)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i1_2_lut_rep_389_3_lut.init = 16'hfdfd;
    LUT4 i1_2_lut_rep_371_3_lut_4_lut (.A(\spi_cmd[1] ), .B(n29141), .C(\spi_cmd[2] ), 
         .D(\spi_addr[0] ), .Z(n29099)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i1_2_lut_rep_371_3_lut_4_lut.init = 16'hfffd;
    LUT4 i14368_3_lut (.A(n19491), .B(resetn_c), .C(n19337), .Z(clk_1MHz_enable_99)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B))) */ ;
    defparam i14368_3_lut.init = 16'h4c4c;
    LUT4 i22619_4_lut (.A(NSL), .B(n19337), .C(n19491), .D(n11859), 
         .Z(NSL_N_4146)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C+(D))))) */ ;
    defparam i22619_4_lut.init = 16'h3b37;
    LUT4 i1_2_lut_rep_375_3_lut_4_lut (.A(\spi_cmd[1] ), .B(n29141), .C(n13489), 
         .D(\spi_addr[0] ), .Z(n29103)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i1_2_lut_rep_375_3_lut_4_lut.init = 16'hfffd;
    LUT4 i1_2_lut_rep_381_3_lut_4_lut (.A(\spi_cmd[1] ), .B(n29141), .C(n18550), 
         .D(\spi_addr[0] ), .Z(n29109)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/s_links/sources/slot_cards/stepper.v(204[15:41])
    defparam i1_2_lut_rep_381_3_lut_4_lut.init = 16'hffdf;
    LUT4 i1_2_lut_adj_478 (.A(Cnt_NSL[7]), .B(Cnt_NSL[8]), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_478.init = 16'heeee;
    LUT4 i2_4_lut_adj_479 (.A(n29253), .B(Cnt[5]), .C(n13386), .D(n19453), 
         .Z(n19423)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i2_4_lut_adj_479.init = 16'hfefa;
    FD1P3IX MA_Temp_474 (.D(MA_Temp_N_3938), .SP(clk_1MHz_enable_378), .CD(n29239), 
            .CK(clk_1MHz), .Q(MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam MA_Temp_474.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \stepper(DEV_ID=4,UART_ADDRESS_WIDTH=4) 
//

module \stepper(DEV_ID=4,UART_ADDRESS_WIDTH=4)  (GND_net, clk_1MHz, clk_1MHz_enable_66, 
            n29239, \SLO_buf[0] , pin_io_out_48, spi_data_out_r_39__N_5174, 
            clk, \spi_data_out_r_39__N_5436[0] , mode_adj_10, clk_enable_359, 
            n29762, n29091, \SLO_buf[13] , \SLO_buf[12] , \SLO_buf[11] , 
            \SLO_buf[10] , \spi_data_out_r_39__N_5436[35] , \spi_data_out_r_39__N_5436[34] , 
            \spi_data_out_r_39__N_5436[33] , \spi_data_out_r_39__N_5436[32] , 
            \spi_data_out_r_39__N_5436[15] , \spi_data_out_r_39__N_5436[14] , 
            \spi_data_out_r_39__N_5436[13] , \spi_data_out_r_39__N_5436[12] , 
            \spi_data_out_r_39__N_5436[11] , \spi_data_out_r_39__N_5436[10] , 
            \spi_data_out_r_39__N_5436[9] , \spi_data_out_r_39__N_5436[8] , 
            \spi_data_out_r_39__N_5436[7] , \spi_data_out_r_39__N_5436[6] , 
            \spi_data_out_r_39__N_5436[5] , \spi_data_out_r_39__N_5436[4] , 
            \spi_data_out_r_39__N_5436[3] , \spi_data_out_r_39__N_5436[2] , 
            \spi_data_out_r_39__N_5436[1] , \SLO_buf[29] , \SLO_buf[28] , 
            \SLO_buf[27] , \SLO_buf[26] , \SLO_buf[25] , \SLO_buf[24] , 
            \SLO_buf[23] , \SLO_buf[22] , \SLO_buf[21] , \SLO_buf[20] , 
            \SLO_buf[19] , \SLO_buf[18] , \SLO_buf[17] , \SLO_buf[16] , 
            \SLO_buf[15] , \SLO_buf[14] , \SLO_buf[9] , \SLO_buf[8] , 
            \SLO_buf[7] , \SLO_buf[6] , \SLO_buf[5] , \SLO_buf[4] , 
            \SLO_buf[3] , \SLO_buf[2] , \SLO_buf[1] , spi_data_out_r_39__N_5214, 
            spi_data_out_r_39__N_5507, digital_output_r, clk_enable_206, 
            \spi_data_r[0] , n29207, n29189, n5, C_5_c_c, n26965, 
            n19381, resetn_c, n29204, OW_ID_N_5482, n29285, mode, 
            n27477, n25411, pin_io_out_49, \quad_b[4] , \quad_a[4] , 
            n1, n1_adj_9, \spi_data_r[1] , \spi_data_r[2] , pin_io_out_44, 
            n29224, quad_homing, n26938, reset_r, clk_enable_526, 
            n29077) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input clk_1MHz;
    input clk_1MHz_enable_66;
    input n29239;
    output \SLO_buf[0] ;
    input pin_io_out_48;
    output [39:0]spi_data_out_r_39__N_5174;
    input clk;
    input \spi_data_out_r_39__N_5436[0] ;
    output [2:0]mode_adj_10;
    input clk_enable_359;
    input n29762;
    input n29091;
    output \SLO_buf[13] ;
    output \SLO_buf[12] ;
    output \SLO_buf[11] ;
    output \SLO_buf[10] ;
    input \spi_data_out_r_39__N_5436[35] ;
    input \spi_data_out_r_39__N_5436[34] ;
    input \spi_data_out_r_39__N_5436[33] ;
    input \spi_data_out_r_39__N_5436[32] ;
    input \spi_data_out_r_39__N_5436[15] ;
    input \spi_data_out_r_39__N_5436[14] ;
    input \spi_data_out_r_39__N_5436[13] ;
    input \spi_data_out_r_39__N_5436[12] ;
    input \spi_data_out_r_39__N_5436[11] ;
    input \spi_data_out_r_39__N_5436[10] ;
    input \spi_data_out_r_39__N_5436[9] ;
    input \spi_data_out_r_39__N_5436[8] ;
    input \spi_data_out_r_39__N_5436[7] ;
    input \spi_data_out_r_39__N_5436[6] ;
    input \spi_data_out_r_39__N_5436[5] ;
    input \spi_data_out_r_39__N_5436[4] ;
    input \spi_data_out_r_39__N_5436[3] ;
    input \spi_data_out_r_39__N_5436[2] ;
    input \spi_data_out_r_39__N_5436[1] ;
    output \SLO_buf[29] ;
    output \SLO_buf[28] ;
    output \SLO_buf[27] ;
    output \SLO_buf[26] ;
    output \SLO_buf[25] ;
    output \SLO_buf[24] ;
    output \SLO_buf[23] ;
    output \SLO_buf[22] ;
    output \SLO_buf[21] ;
    output \SLO_buf[20] ;
    output \SLO_buf[19] ;
    output \SLO_buf[18] ;
    output \SLO_buf[17] ;
    output \SLO_buf[16] ;
    output \SLO_buf[15] ;
    output \SLO_buf[14] ;
    output \SLO_buf[9] ;
    output \SLO_buf[8] ;
    output \SLO_buf[7] ;
    output \SLO_buf[6] ;
    output \SLO_buf[5] ;
    output \SLO_buf[4] ;
    output \SLO_buf[3] ;
    output \SLO_buf[2] ;
    output \SLO_buf[1] ;
    output spi_data_out_r_39__N_5214;
    input spi_data_out_r_39__N_5507;
    output digital_output_r;
    input clk_enable_206;
    input \spi_data_r[0] ;
    output n29207;
    input n29189;
    input n5;
    input C_5_c_c;
    output n26965;
    output n19381;
    input resetn_c;
    input n29204;
    output OW_ID_N_5482;
    input n29285;
    input mode;
    output n27477;
    output n25411;
    input pin_io_out_49;
    output \quad_b[4] ;
    output \quad_a[4] ;
    output n1;
    output n1_adj_9;
    input \spi_data_r[1] ;
    input \spi_data_r[2] ;
    input pin_io_out_44;
    input n29224;
    input [1:0]quad_homing;
    output n26938;
    output reset_r;
    input clk_enable_526;
    input n29077;
    
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire MA_Temp_N_5291 /* synthesis is_inv_clock=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    wire clk_1MHz_derived_134 /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz_derived_134 */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire MA_Temp /* synthesis is_clock=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(57[5:12])
    
    wire n25021;
    wire [11:0]Cnt_NSL;   // c:/s_links/sources/slot_cards/stepper.v(61[12:19])
    wire [11:0]n1290;
    
    wire n25022;
    wire [51:0]SLO;   // c:/s_links/sources/slot_cards/stepper.v(63[12:15])
    
    wire clk_1MHz_derived_134_enable_46;
    wire [7:0]Cnt;   // c:/s_links/sources/slot_cards/stepper.v(62[11:14])
    
    wire clk_1MHz_enable_349;
    wire [7:0]n199;
    wire [51:0]SLO_buf;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire clk_1MHz_derived_134_enable_27, n29140, n25020, n25019, n19433, 
        n19525;
    wire [31:0]n153;
    
    wire n28931, n28928, n29206, MA_Temp_N_5294, n29281, n28929, 
        n4, clk_1MHz_enable_341, n29164, n13384, n27462, n25018, 
        n25017, n25016, n25015, clk_1MHz_enable_214, NSL, n11805, 
        NSL_N_5502, n28930, n29289, n29290, n19461, n25024, n25023;
    
    CCU2D add_551_7 (.A0(Cnt_NSL[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25021), .COUT(n25022), .S0(n1290[5]), .S1(n1290[6]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_7.INIT0 = 16'h5aaa;
    defparam add_551_7.INIT1 = 16'h5aaa;
    defparam add_551_7.INJECT1_0 = "NO";
    defparam add_551_7.INJECT1_1 = "NO";
    FD1P3IX Cnt_NSL__i0 (.D(n1290[0]), .SP(clk_1MHz_enable_66), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i0.GSR = "DISABLED";
    FD1S3AX SLO_buf_i1 (.D(SLO[0]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i1.GSR = "DISABLED";
    FD1P3AX SLO_i0 (.D(pin_io_out_48), .SP(clk_1MHz_derived_134_enable_46), 
            .CK(clk_1MHz_derived_134), .Q(SLO[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i0 (.D(\spi_data_out_r_39__N_5436[0] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i0.GSR = "DISABLED";
    FD1P3IX mode__i0 (.D(n29762), .SP(clk_enable_359), .CD(n29239), .CK(clk), 
            .Q(mode_adj_10[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i0.GSR = "DISABLED";
    FD1P3IX Cnt__i0 (.D(n199[0]), .SP(clk_1MHz_enable_349), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i0.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i39 (.D(\SLO_buf[13] ), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i39.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i38 (.D(\SLO_buf[12] ), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i38.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i37 (.D(\SLO_buf[11] ), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i37.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i36 (.D(\SLO_buf[10] ), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i36.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i35 (.D(\spi_data_out_r_39__N_5436[35] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i35.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i34 (.D(\spi_data_out_r_39__N_5436[34] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i34.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i33 (.D(\spi_data_out_r_39__N_5436[33] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i33.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_5436[32] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i31 (.D(SLO_buf[45]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i30 (.D(SLO_buf[44]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i29 (.D(SLO_buf[43]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i28 (.D(SLO_buf[42]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i27 (.D(SLO_buf[41]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i26 (.D(SLO_buf[40]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i25 (.D(SLO_buf[39]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i24 (.D(SLO_buf[38]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i23 (.D(SLO_buf[37]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i22 (.D(SLO_buf[36]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i21 (.D(SLO_buf[35]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i20 (.D(SLO_buf[34]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i19 (.D(SLO_buf[33]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i18 (.D(SLO_buf[32]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i17 (.D(SLO_buf[31]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i16 (.D(SLO_buf[30]), .CK(clk), .CD(n29091), 
            .Q(spi_data_out_r_39__N_5174[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_5436[15] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_5436[14] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_5436[13] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_5436[12] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_5436[11] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_5436[10] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_5436[9] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_5436[8] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_5436[7] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_5436[6] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_5436[5] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_5436[4] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_5436[3] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_5436[2] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_5436[1] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5174[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1P3IX SLO_i45 (.D(SLO[44]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i45.GSR = "DISABLED";
    FD1P3IX SLO_i44 (.D(SLO[43]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i44.GSR = "DISABLED";
    FD1P3IX SLO_i43 (.D(SLO[42]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i43.GSR = "DISABLED";
    FD1P3IX SLO_i42 (.D(SLO[41]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i42.GSR = "DISABLED";
    FD1P3IX SLO_i41 (.D(SLO[40]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i41.GSR = "DISABLED";
    FD1P3IX SLO_i40 (.D(SLO[39]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i40.GSR = "DISABLED";
    FD1P3IX SLO_i39 (.D(SLO[38]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i39.GSR = "DISABLED";
    FD1P3IX SLO_i38 (.D(SLO[37]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i38.GSR = "DISABLED";
    FD1P3IX SLO_i37 (.D(SLO[36]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i37.GSR = "DISABLED";
    FD1P3IX SLO_i36 (.D(SLO[35]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i36.GSR = "DISABLED";
    FD1P3IX SLO_i35 (.D(SLO[34]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i35.GSR = "DISABLED";
    FD1P3IX SLO_i34 (.D(SLO[33]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i34.GSR = "DISABLED";
    FD1P3IX SLO_i33 (.D(SLO[32]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i33.GSR = "DISABLED";
    FD1P3IX SLO_i32 (.D(SLO[31]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i32.GSR = "DISABLED";
    FD1P3IX SLO_i31 (.D(SLO[30]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i31.GSR = "DISABLED";
    FD1P3IX SLO_i30 (.D(SLO[29]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i30.GSR = "DISABLED";
    FD1P3IX SLO_i29 (.D(SLO[28]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i29.GSR = "DISABLED";
    FD1P3IX SLO_i28 (.D(SLO[27]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i28.GSR = "DISABLED";
    FD1P3IX SLO_i27 (.D(SLO[26]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i27.GSR = "DISABLED";
    FD1P3IX SLO_i26 (.D(SLO[25]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i26.GSR = "DISABLED";
    FD1P3IX SLO_i25 (.D(SLO[24]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i25.GSR = "DISABLED";
    FD1P3IX SLO_i24 (.D(SLO[23]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i24.GSR = "DISABLED";
    FD1P3IX SLO_i23 (.D(SLO[22]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i23.GSR = "DISABLED";
    FD1P3IX SLO_i22 (.D(SLO[21]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i22.GSR = "DISABLED";
    FD1P3IX SLO_i21 (.D(SLO[20]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i21.GSR = "DISABLED";
    FD1P3IX SLO_i20 (.D(SLO[19]), .SP(clk_1MHz_derived_134_enable_27), .CD(n29140), 
            .CK(clk_1MHz_derived_134), .Q(SLO[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i20.GSR = "DISABLED";
    FD1P3AX SLO_i19 (.D(SLO[18]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i19.GSR = "DISABLED";
    FD1P3AX SLO_i18 (.D(SLO[17]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i18.GSR = "DISABLED";
    FD1P3AX SLO_i17 (.D(SLO[16]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i17.GSR = "DISABLED";
    FD1P3AX SLO_i16 (.D(SLO[15]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i16.GSR = "DISABLED";
    FD1P3AX SLO_i15 (.D(SLO[14]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i15.GSR = "DISABLED";
    FD1P3AX SLO_i14 (.D(SLO[13]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i14.GSR = "DISABLED";
    FD1P3AX SLO_i13 (.D(SLO[12]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i13.GSR = "DISABLED";
    FD1P3AX SLO_i12 (.D(SLO[11]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i12.GSR = "DISABLED";
    FD1P3AX SLO_i11 (.D(SLO[10]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i11.GSR = "DISABLED";
    FD1P3AX SLO_i10 (.D(SLO[9]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i10.GSR = "DISABLED";
    FD1P3AX SLO_i9 (.D(SLO[8]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i9.GSR = "DISABLED";
    FD1P3AX SLO_i8 (.D(SLO[7]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i8.GSR = "DISABLED";
    FD1P3AX SLO_i7 (.D(SLO[6]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i7.GSR = "DISABLED";
    FD1P3AX SLO_i6 (.D(SLO[5]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i6.GSR = "DISABLED";
    FD1P3AX SLO_i5 (.D(SLO[4]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i5.GSR = "DISABLED";
    FD1P3AX SLO_i4 (.D(SLO[3]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i4.GSR = "DISABLED";
    FD1P3AX SLO_i3 (.D(SLO[2]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i3.GSR = "DISABLED";
    FD1P3AX SLO_i2 (.D(SLO[1]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i2.GSR = "DISABLED";
    FD1P3AX SLO_i1 (.D(SLO[0]), .SP(clk_1MHz_derived_134_enable_46), .CK(clk_1MHz_derived_134), 
            .Q(SLO[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i1.GSR = "DISABLED";
    FD1S3AX SLO_buf_i46 (.D(SLO[45]), .CK(MA_Temp_N_5291), .Q(SLO_buf[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i46.GSR = "DISABLED";
    FD1S3AX SLO_buf_i45 (.D(SLO[44]), .CK(MA_Temp_N_5291), .Q(SLO_buf[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i45.GSR = "DISABLED";
    FD1S3AX SLO_buf_i44 (.D(SLO[43]), .CK(MA_Temp_N_5291), .Q(SLO_buf[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i44.GSR = "DISABLED";
    FD1S3AX SLO_buf_i43 (.D(SLO[42]), .CK(MA_Temp_N_5291), .Q(SLO_buf[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i43.GSR = "DISABLED";
    FD1S3AX SLO_buf_i42 (.D(SLO[41]), .CK(MA_Temp_N_5291), .Q(SLO_buf[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i42.GSR = "DISABLED";
    FD1S3AX SLO_buf_i41 (.D(SLO[40]), .CK(MA_Temp_N_5291), .Q(SLO_buf[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i41.GSR = "DISABLED";
    FD1S3AX SLO_buf_i40 (.D(SLO[39]), .CK(MA_Temp_N_5291), .Q(SLO_buf[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i40.GSR = "DISABLED";
    FD1S3AX SLO_buf_i39 (.D(SLO[38]), .CK(MA_Temp_N_5291), .Q(SLO_buf[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i39.GSR = "DISABLED";
    FD1S3AX SLO_buf_i38 (.D(SLO[37]), .CK(MA_Temp_N_5291), .Q(SLO_buf[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i38.GSR = "DISABLED";
    FD1S3AX SLO_buf_i37 (.D(SLO[36]), .CK(MA_Temp_N_5291), .Q(SLO_buf[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i37.GSR = "DISABLED";
    FD1S3AX SLO_buf_i36 (.D(SLO[35]), .CK(MA_Temp_N_5291), .Q(SLO_buf[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i36.GSR = "DISABLED";
    FD1S3AX SLO_buf_i35 (.D(SLO[34]), .CK(MA_Temp_N_5291), .Q(SLO_buf[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i35.GSR = "DISABLED";
    FD1S3AX SLO_buf_i34 (.D(SLO[33]), .CK(MA_Temp_N_5291), .Q(SLO_buf[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i34.GSR = "DISABLED";
    FD1S3AX SLO_buf_i33 (.D(SLO[32]), .CK(MA_Temp_N_5291), .Q(SLO_buf[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i33.GSR = "DISABLED";
    FD1S3AX SLO_buf_i32 (.D(SLO[31]), .CK(MA_Temp_N_5291), .Q(SLO_buf[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i32.GSR = "DISABLED";
    FD1S3AX SLO_buf_i31 (.D(SLO[30]), .CK(MA_Temp_N_5291), .Q(SLO_buf[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i31.GSR = "DISABLED";
    FD1S3AX SLO_buf_i30 (.D(SLO[29]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i30.GSR = "DISABLED";
    FD1S3AX SLO_buf_i29 (.D(SLO[28]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i29.GSR = "DISABLED";
    FD1S3AX SLO_buf_i28 (.D(SLO[27]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i28.GSR = "DISABLED";
    FD1S3AX SLO_buf_i27 (.D(SLO[26]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i27.GSR = "DISABLED";
    FD1S3AX SLO_buf_i26 (.D(SLO[25]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i26.GSR = "DISABLED";
    FD1S3AX SLO_buf_i25 (.D(SLO[24]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i25.GSR = "DISABLED";
    FD1S3AX SLO_buf_i24 (.D(SLO[23]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i24.GSR = "DISABLED";
    FD1S3AX SLO_buf_i23 (.D(SLO[22]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i23.GSR = "DISABLED";
    FD1S3AX SLO_buf_i22 (.D(SLO[21]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i22.GSR = "DISABLED";
    FD1S3AX SLO_buf_i21 (.D(SLO[20]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i21.GSR = "DISABLED";
    FD1S3AX SLO_buf_i20 (.D(SLO[19]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i20.GSR = "DISABLED";
    FD1S3AX SLO_buf_i19 (.D(SLO[18]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i19.GSR = "DISABLED";
    FD1S3AX SLO_buf_i18 (.D(SLO[17]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i18.GSR = "DISABLED";
    FD1S3AX SLO_buf_i17 (.D(SLO[16]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i17.GSR = "DISABLED";
    FD1S3AX SLO_buf_i16 (.D(SLO[15]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i16.GSR = "DISABLED";
    FD1S3AX SLO_buf_i15 (.D(SLO[14]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i15.GSR = "DISABLED";
    FD1S3AX SLO_buf_i14 (.D(SLO[13]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i14.GSR = "DISABLED";
    FD1S3AX SLO_buf_i13 (.D(SLO[12]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i13.GSR = "DISABLED";
    FD1S3AX SLO_buf_i12 (.D(SLO[11]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i12.GSR = "DISABLED";
    FD1S3AX SLO_buf_i11 (.D(SLO[10]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i11.GSR = "DISABLED";
    FD1S3AX SLO_buf_i10 (.D(SLO[9]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i10.GSR = "DISABLED";
    FD1S3AX SLO_buf_i9 (.D(SLO[8]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i9.GSR = "DISABLED";
    FD1S3AX SLO_buf_i8 (.D(SLO[7]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i8.GSR = "DISABLED";
    FD1S3AX SLO_buf_i7 (.D(SLO[6]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i7.GSR = "DISABLED";
    FD1S3AX SLO_buf_i6 (.D(SLO[5]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i6.GSR = "DISABLED";
    FD1S3AX SLO_buf_i5 (.D(SLO[4]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i5.GSR = "DISABLED";
    FD1S3AX SLO_buf_i4 (.D(SLO[3]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i4.GSR = "DISABLED";
    FD1S3AX SLO_buf_i3 (.D(SLO[2]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i3.GSR = "DISABLED";
    FD1S3AX SLO_buf_i2 (.D(SLO[1]), .CK(MA_Temp_N_5291), .Q(\SLO_buf[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i2.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i11 (.D(n1290[11]), .SP(clk_1MHz_enable_66), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i11.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i10 (.D(n1290[10]), .SP(clk_1MHz_enable_66), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i10.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i9 (.D(n1290[9]), .SP(clk_1MHz_enable_66), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i9.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i8 (.D(n1290[8]), .SP(clk_1MHz_enable_66), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i8.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i7 (.D(n1290[7]), .SP(clk_1MHz_enable_66), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i7.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i6 (.D(n1290[6]), .SP(clk_1MHz_enable_66), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i6.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i5 (.D(n1290[5]), .SP(clk_1MHz_enable_66), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i5.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i4 (.D(n1290[4]), .SP(clk_1MHz_enable_66), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i4.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i3 (.D(n1290[3]), .SP(clk_1MHz_enable_66), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i3.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i2 (.D(n1290[2]), .SP(clk_1MHz_enable_66), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i2.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i1 (.D(n1290[1]), .SP(clk_1MHz_enable_66), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i1.GSR = "DISABLED";
    CCU2D add_551_5 (.A0(Cnt_NSL[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25020), .COUT(n25021), .S0(n1290[3]), .S1(n1290[4]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_5.INIT0 = 16'h5aaa;
    defparam add_551_5.INIT1 = 16'h5aaa;
    defparam add_551_5.INJECT1_0 = "NO";
    defparam add_551_5.INJECT1_1 = "NO";
    CCU2D add_551_3 (.A0(Cnt_NSL[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25019), .COUT(n25020), .S0(n1290[1]), .S1(n1290[2]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_3.INIT0 = 16'h5aaa;
    defparam add_551_3.INIT1 = 16'h5aaa;
    defparam add_551_3.INJECT1_0 = "NO";
    defparam add_551_3.INJECT1_1 = "NO";
    LUT4 i13665_2_lut_3_lut (.A(n19433), .B(n19525), .C(n153[0]), .Z(n199[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13665_2_lut_3_lut.init = 16'h7070;
    LUT4 i13734_2_lut_3_lut (.A(n19433), .B(n19525), .C(n153[1]), .Z(n199[1])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13734_2_lut_3_lut.init = 16'h7070;
    LUT4 i13733_2_lut_3_lut (.A(n19433), .B(n19525), .C(n153[2]), .Z(n199[2])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13733_2_lut_3_lut.init = 16'h7070;
    LUT4 n28931_bdd_3_lut (.A(n28931), .B(n28928), .C(n29206), .Z(MA_Temp_N_5294)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28931_bdd_3_lut.init = 16'hcaca;
    LUT4 i13732_2_lut_3_lut (.A(n19433), .B(n19525), .C(n153[3]), .Z(n199[3])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13732_2_lut_3_lut.init = 16'h7070;
    LUT4 i13731_2_lut_3_lut (.A(n19433), .B(n19525), .C(n153[4]), .Z(n199[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13731_2_lut_3_lut.init = 16'h7070;
    LUT4 i13730_2_lut_3_lut (.A(n19433), .B(n19525), .C(n153[5]), .Z(n199[5])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13730_2_lut_3_lut.init = 16'h7070;
    FD1S3IX i159_483 (.D(spi_data_out_r_39__N_5507), .CK(clk), .CD(n29239), 
            .Q(spi_data_out_r_39__N_5214)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam i159_483.GSR = "DISABLED";
    LUT4 i13729_2_lut_3_lut (.A(n19433), .B(n19525), .C(n153[6]), .Z(n199[6])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13729_2_lut_3_lut.init = 16'h7070;
    LUT4 i13728_2_lut_3_lut (.A(n19433), .B(n19525), .C(n153[7]), .Z(n199[7])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13728_2_lut_3_lut.init = 16'h7070;
    LUT4 n19433_bdd_4_lut_23359 (.A(n19433), .B(n29281), .C(MA_Temp), 
         .D(Cnt[5]), .Z(n28929)) /* synthesis lut_function=(!(A+(B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam n19433_bdd_4_lut_23359.init = 16'h1450;
    LUT4 n19433_bdd_3_lut_23111 (.A(n19433), .B(n19525), .C(MA_Temp), 
         .Z(n28928)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam n19433_bdd_3_lut_23111.init = 16'h7070;
    FD1P3IX digital_output_r_481 (.D(\spi_data_r[0] ), .SP(clk_enable_206), 
            .CD(n29239), .CK(clk), .Q(digital_output_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam digital_output_r_481.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut (.A(n29207), .B(n29189), .C(n5), .D(C_5_c_c), 
         .Z(n26965)) /* synthesis lut_function=((B (C+(D))+!B (C))+!A) */ ;   // c:/s_links/sources/slot_cards/stepper.v(71[15:39])
    defparam i1_4_lut_4_lut.init = 16'hfdf5;
    LUT4 i2_4_lut (.A(Cnt_NSL[11]), .B(Cnt_NSL[9]), .C(Cnt_NSL[10]), .D(n4), 
         .Z(n19381)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'ha080;
    LUT4 i1_2_lut (.A(Cnt_NSL[7]), .B(Cnt_NSL[8]), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i22773_2_lut_rep_424 (.A(n19381), .B(resetn_c), .Z(clk_1MHz_enable_349)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i22773_2_lut_rep_424.init = 16'hbbbb;
    LUT4 i22878_2_lut_2_lut_3_lut_4_lut (.A(n19381), .B(resetn_c), .C(n19525), 
         .D(n19433), .Z(clk_1MHz_enable_341)) /* synthesis lut_function=(!(A (C (D))+!A (B+(C (D))))) */ ;
    defparam i22878_2_lut_2_lut_3_lut_4_lut.init = 16'h0bbb;
    LUT4 i117_4_lut (.A(n29164), .B(n13384), .C(Cnt[1]), .D(Cnt[4]), 
         .Z(clk_1MHz_derived_134_enable_27)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(132[15:49])
    defparam i117_4_lut.init = 16'h3332;
    LUT4 i1_2_lut_adj_371 (.A(Cnt[2]), .B(Cnt[3]), .Z(n27462)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_adj_371.init = 16'heeee;
    LUT4 i1_4_lut (.A(n29204), .B(OW_ID_N_5482), .C(n29285), .D(mode), 
         .Z(n27477)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(94[6:59])
    defparam i1_4_lut.init = 16'h5554;
    CCU2D add_551_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n25019), .S1(n1290[0]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_1.INIT0 = 16'hF000;
    defparam add_551_1.INIT1 = 16'h5555;
    defparam add_551_1.INJECT1_0 = "NO";
    defparam add_551_1.INJECT1_1 = "NO";
    CCU2D add_552_9 (.A0(Cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25018), 
          .S0(n153[7]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_9.INIT0 = 16'h5aaa;
    defparam add_552_9.INIT1 = 16'h0000;
    defparam add_552_9.INJECT1_0 = "NO";
    defparam add_552_9.INJECT1_1 = "NO";
    CCU2D add_552_7 (.A0(Cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25017), 
          .COUT(n25018), .S0(n153[5]), .S1(n153[6]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_7.INIT0 = 16'h5aaa;
    defparam add_552_7.INIT1 = 16'h5aaa;
    defparam add_552_7.INJECT1_0 = "NO";
    defparam add_552_7.INJECT1_1 = "NO";
    CCU2D add_552_5 (.A0(Cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25016), 
          .COUT(n25017), .S0(n153[3]), .S1(n153[4]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_5.INIT0 = 16'h5aaa;
    defparam add_552_5.INIT1 = 16'h5aaa;
    defparam add_552_5.INJECT1_0 = "NO";
    defparam add_552_5.INJECT1_1 = "NO";
    CCU2D add_552_3 (.A0(Cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25015), 
          .COUT(n25016), .S0(n153[1]), .S1(n153[2]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_3.INIT0 = 16'h5aaa;
    defparam add_552_3.INIT1 = 16'h5aaa;
    defparam add_552_3.INJECT1_0 = "NO";
    defparam add_552_3.INJECT1_1 = "NO";
    CCU2D add_552_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n25015), 
          .S1(n153[0]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_1.INIT0 = 16'hF000;
    defparam add_552_1.INIT1 = 16'h5555;
    defparam add_552_1.INJECT1_0 = "NO";
    defparam add_552_1.INJECT1_1 = "NO";
    LUT4 i14372_3_lut (.A(n19525), .B(resetn_c), .C(n19381), .Z(clk_1MHz_enable_214)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B))) */ ;
    defparam i14372_3_lut.init = 16'h4c4c;
    LUT4 i22653_4_lut (.A(NSL), .B(n19381), .C(n19525), .D(n11805), 
         .Z(NSL_N_5502)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C+(D))))) */ ;
    defparam i22653_4_lut.init = 16'h3b37;
    LUT4 i14326_2_lut_rep_553 (.A(Cnt[4]), .B(Cnt[1]), .Z(n29281)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14326_2_lut_rep_553.init = 16'h8888;
    LUT4 n19433_bdd_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(Cnt[5]), .D(MA_Temp), 
         .Z(n28930)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;
    defparam n19433_bdd_3_lut_4_lut.init = 16'hf708;
    LUT4 i1_2_lut_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(n29206), .D(Cnt[5]), 
         .Z(n11805)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut_rep_436_4_lut (.A(n27462), .B(Cnt[0]), .C(n29289), .D(Cnt[5]), 
         .Z(n29164)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_rep_436_4_lut.init = 16'hfffe;
    LUT4 i22820_3_lut_3_lut_3_lut_4_lut (.A(mode_adj_10[0]), .B(n29290), 
         .C(n29285), .D(n29189), .Z(n25411)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i22820_3_lut_3_lut_3_lut_4_lut.init = 16'h000d;
    FD1P3AX NSL_476 (.D(NSL_N_5502), .SP(clk_1MHz_enable_214), .CK(clk_1MHz), 
            .Q(NSL)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam NSL_476.GSR = "DISABLED";
    LUT4 i2_4_lut_adj_372 (.A(n29289), .B(Cnt[5]), .C(n13384), .D(n19461), 
         .Z(n19433)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i2_4_lut_adj_372.init = 16'hfefa;
    LUT4 Select_4096_i1_2_lut_3_lut_4_lut (.A(mode_adj_10[0]), .B(mode_adj_10[2]), 
         .C(pin_io_out_49), .D(mode_adj_10[1]), .Z(\quad_b[4] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam Select_4096_i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 Select_4089_i1_2_lut_3_lut_4_lut (.A(mode_adj_10[0]), .B(mode_adj_10[2]), 
         .C(pin_io_out_48), .D(mode_adj_10[1]), .Z(\quad_a[4] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam Select_4089_i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_3_lut (.A(mode_adj_10[0]), .B(mode_adj_10[2]), .C(mode_adj_10[1]), 
         .Z(OW_ID_N_5482)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_561 (.A(Cnt[6]), .B(Cnt[7]), .Z(n29289)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_rep_561.init = 16'heeee;
    LUT4 i2_3_lut_rep_478_4_lut (.A(Cnt[6]), .B(Cnt[7]), .C(Cnt[0]), .D(n27462), 
         .Z(n29206)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i2_3_lut_rep_478_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_562 (.A(mode_adj_10[1]), .B(mode_adj_10[2]), .Z(n29290)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_rep_562.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_479_3_lut (.A(mode_adj_10[1]), .B(mode_adj_10[2]), 
         .C(mode_adj_10[0]), .Z(n29207)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_rep_479_3_lut.init = 16'hbfbf;
    LUT4 Select_3906_i1_2_lut_2_lut_3_lut_4_lut (.A(mode_adj_10[1]), .B(mode_adj_10[2]), 
         .C(NSL), .D(mode_adj_10[0]), .Z(n1)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam Select_3906_i1_2_lut_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_3_lut_adj_373 (.A(mode_adj_10[1]), .B(mode_adj_10[2]), 
         .C(mode_adj_10[0]), .Z(n13384)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_3_lut_adj_373.init = 16'hfbfb;
    LUT4 equal_139_i6_1_lut_rep_412_2_lut_3_lut (.A(mode_adj_10[1]), .B(mode_adj_10[2]), 
         .C(mode_adj_10[0]), .Z(n29140)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam equal_139_i6_1_lut_rep_412_2_lut_3_lut.init = 16'h4040;
    LUT4 i5013_2_lut_3_lut_4_lut (.A(mode_adj_10[1]), .B(mode_adj_10[2]), 
         .C(clk_1MHz_derived_134_enable_27), .D(mode_adj_10[0]), .Z(clk_1MHz_derived_134_enable_46)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i5013_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i22656_2_lut_rep_566 (.A(MA_Temp), .B(clk_1MHz), .Z(clk_1MHz_derived_134)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[13:34])
    defparam i22656_2_lut_rep_566.init = 16'h7777;
    LUT4 Select_3903_i1_2_lut_3_lut (.A(MA_Temp), .B(clk_1MHz), .C(mode_adj_10[2]), 
         .Z(n1_adj_9)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[13:34])
    defparam Select_3903_i1_2_lut_3_lut.init = 16'h7070;
    LUT4 i3_4_lut (.A(n19461), .B(Cnt[5]), .C(n29207), .D(n29289), .Z(n19525)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i14521_4_lut (.A(Cnt[0]), .B(Cnt[4]), .C(n27462), .D(Cnt[1]), 
         .Z(n19461)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i14521_4_lut.init = 16'hc8c0;
    FD1P3IX MA_Temp_474 (.D(MA_Temp_N_5294), .SP(clk_1MHz_enable_341), .CD(n29239), 
            .CK(clk_1MHz), .Q(MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam MA_Temp_474.GSR = "DISABLED";
    FD1P3IX mode__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_359), .CD(n29239), 
            .CK(clk), .Q(mode_adj_10[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i1.GSR = "DISABLED";
    FD1P3IX mode__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_359), .CD(n29239), 
            .CK(clk), .Q(mode_adj_10[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i1 (.D(n199[1]), .SP(clk_1MHz_enable_349), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i1.GSR = "DISABLED";
    FD1P3IX Cnt__i2 (.D(n199[2]), .SP(clk_1MHz_enable_349), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i3 (.D(n199[3]), .SP(clk_1MHz_enable_349), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i3.GSR = "DISABLED";
    FD1P3IX Cnt__i4 (.D(n199[4]), .SP(clk_1MHz_enable_349), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i4.GSR = "DISABLED";
    FD1P3IX Cnt__i5 (.D(n199[5]), .SP(clk_1MHz_enable_349), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i5.GSR = "DISABLED";
    FD1P3IX Cnt__i6 (.D(n199[6]), .SP(clk_1MHz_enable_349), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i6.GSR = "DISABLED";
    FD1P3IX Cnt__i7 (.D(n199[7]), .SP(clk_1MHz_enable_349), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i7.GSR = "DISABLED";
    CCU2D add_551_13 (.A0(Cnt_NSL[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25024), 
          .S0(n1290[11]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_13.INIT0 = 16'h5aaa;
    defparam add_551_13.INIT1 = 16'h0000;
    defparam add_551_13.INJECT1_0 = "NO";
    defparam add_551_13.INJECT1_1 = "NO";
    CCU2D add_551_11 (.A0(Cnt_NSL[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25023), .COUT(n25024), .S0(n1290[9]), .S1(n1290[10]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_11.INIT0 = 16'h5aaa;
    defparam add_551_11.INIT1 = 16'h5aaa;
    defparam add_551_11.INJECT1_0 = "NO";
    defparam add_551_11.INJECT1_1 = "NO";
    CCU2D add_551_9 (.A0(Cnt_NSL[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25022), .COUT(n25023), .S0(n1290[7]), .S1(n1290[8]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_9.INIT0 = 16'h5aaa;
    defparam add_551_9.INIT1 = 16'h5aaa;
    defparam add_551_9.INJECT1_0 = "NO";
    defparam add_551_9.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_374 (.A(pin_io_out_44), .B(n29224), .C(quad_homing[1]), 
         .D(quad_homing[0]), .Z(n26938)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(75[8:17])
    defparam i1_4_lut_adj_374.init = 16'h0200;
    INV i23372 (.A(MA_Temp), .Z(MA_Temp_N_5291));
    FD1P3IX reset_r_480 (.D(n29077), .SP(clk_enable_526), .CD(n29239), 
            .CK(clk), .Q(reset_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam reset_r_480.GSR = "DISABLED";
    PFUMX i23112 (.BLUT(n28930), .ALUT(n28929), .C0(n19525), .Z(n28931));
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \rs232(DEV_ID=4,UART_ADDRESS_WIDTH=4) 
//

module \rs232(DEV_ID=4,UART_ADDRESS_WIDTH=4)  (\spi_addr_r[0] , \spi_cmd_r[1] , 
            n29255, n29256, n65, n29083, clk, clk_enable_200, n29239, 
            \spi_data_r[0] , C_3_c_2, n29282, C_4_c_3, n29189) /* synthesis syn_module_defined=1 */ ;
    input \spi_addr_r[0] ;
    input \spi_cmd_r[1] ;
    output n29255;
    input n29256;
    input n65;
    output n29083;
    input clk;
    input clk_enable_200;
    input n29239;
    input \spi_data_r[0] ;
    input C_3_c_2;
    input n29282;
    input C_4_c_3;
    output n29189;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    wire mode;
    
    LUT4 i13854_2_lut_rep_527 (.A(\spi_addr_r[0] ), .B(\spi_cmd_r[1] ), 
         .Z(n29255)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i13854_2_lut_rep_527.init = 16'heeee;
    LUT4 i1_2_lut_rep_355_3_lut_4_lut (.A(\spi_addr_r[0] ), .B(\spi_cmd_r[1] ), 
         .C(n29256), .D(n65), .Z(n29083)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_2_lut_rep_355_3_lut_4_lut.init = 16'h1000;
    FD1P3IX mode_26 (.D(\spi_data_r[0] ), .SP(clk_enable_200), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=552, LSE_RLINE=572 */ ;   // c:/s_links/sources/rs232.v(39[8] 47[4])
    defparam mode_26.GSR = "DISABLED";
    LUT4 i2_4_lut_rep_461 (.A(mode), .B(C_3_c_2), .C(n29282), .D(C_4_c_3), 
         .Z(n29189)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2_4_lut_rep_461.init = 16'h0008;
    
endmodule
//
// Verilog Description of module \stepper(DEV_ID=1,UART_ADDRESS_WIDTH=4) 
//

module \stepper(DEV_ID=1,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_30, 
            n29239, \spi_data_r[2] , \spi_data_r[1] , digital_output_r, 
            clk_enable_20, \spi_data_r[0] , spi_data_out_r_39__N_4157, 
            n29094, \SLO_buf[13] , \SLO_buf[12] , \SLO_buf[11] , \SLO_buf[10] , 
            \spi_data_out_r_39__N_4419[35] , \spi_data_out_r_39__N_4419[34] , 
            \spi_data_out_r_39__N_4419[33] , \spi_data_out_r_39__N_4419[32] , 
            \spi_data_out_r_39__N_4419[15] , \spi_data_out_r_39__N_4419[14] , 
            \spi_data_out_r_39__N_4419[13] , \spi_data_out_r_39__N_4419[12] , 
            \spi_data_out_r_39__N_4419[11] , \spi_data_out_r_39__N_4419[10] , 
            \spi_data_out_r_39__N_4419[9] , \spi_data_out_r_39__N_4419[8] , 
            \spi_data_out_r_39__N_4419[7] , \spi_data_out_r_39__N_4419[6] , 
            \spi_data_out_r_39__N_4419[5] , \spi_data_out_r_39__N_4419[4] , 
            \spi_data_out_r_39__N_4419[3] , \spi_data_out_r_39__N_4419[2] , 
            \spi_data_out_r_39__N_4419[1] , pin_io_out_19, \quad_b[1] , 
            pin_io_out_18, \quad_a[1] , GND_net, clk_1MHz, clk_1MHz_enable_91, 
            \SLO_buf[0] , \spi_data_out_r_39__N_4419[0] , spi_data_out_r_39__N_4197, 
            spi_data_out_r_39__N_4490, n29762, \SLO_buf[29] , \SLO_buf[28] , 
            \SLO_buf[27] , \SLO_buf[26] , \SLO_buf[25] , \SLO_buf[24] , 
            \SLO_buf[23] , \SLO_buf[22] , \SLO_buf[21] , \SLO_buf[20] , 
            \SLO_buf[19] , \SLO_buf[18] , \SLO_buf[17] , \SLO_buf[16] , 
            \SLO_buf[15] , \SLO_buf[14] , \SLO_buf[9] , \SLO_buf[8] , 
            \SLO_buf[7] , \SLO_buf[6] , \SLO_buf[5] , \SLO_buf[4] , 
            \SLO_buf[3] , \SLO_buf[2] , \SLO_buf[1] , n19351, resetn_c, 
            n29217, n29315, \cs_decoded[2] , n29306, n8796, OW_ID_N_4464, 
            C_5_c_c, OW_ID_N_4462, reset_r, clk_enable_307, n29097, 
            n1, n1_adj_8) /* synthesis syn_module_defined=1 */ ;
    output [2:0]mode;
    input clk;
    input clk_enable_30;
    input n29239;
    input \spi_data_r[2] ;
    input \spi_data_r[1] ;
    output digital_output_r;
    input clk_enable_20;
    input \spi_data_r[0] ;
    output [39:0]spi_data_out_r_39__N_4157;
    input n29094;
    output \SLO_buf[13] ;
    output \SLO_buf[12] ;
    output \SLO_buf[11] ;
    output \SLO_buf[10] ;
    input \spi_data_out_r_39__N_4419[35] ;
    input \spi_data_out_r_39__N_4419[34] ;
    input \spi_data_out_r_39__N_4419[33] ;
    input \spi_data_out_r_39__N_4419[32] ;
    input \spi_data_out_r_39__N_4419[15] ;
    input \spi_data_out_r_39__N_4419[14] ;
    input \spi_data_out_r_39__N_4419[13] ;
    input \spi_data_out_r_39__N_4419[12] ;
    input \spi_data_out_r_39__N_4419[11] ;
    input \spi_data_out_r_39__N_4419[10] ;
    input \spi_data_out_r_39__N_4419[9] ;
    input \spi_data_out_r_39__N_4419[8] ;
    input \spi_data_out_r_39__N_4419[7] ;
    input \spi_data_out_r_39__N_4419[6] ;
    input \spi_data_out_r_39__N_4419[5] ;
    input \spi_data_out_r_39__N_4419[4] ;
    input \spi_data_out_r_39__N_4419[3] ;
    input \spi_data_out_r_39__N_4419[2] ;
    input \spi_data_out_r_39__N_4419[1] ;
    input pin_io_out_19;
    output \quad_b[1] ;
    input pin_io_out_18;
    output \quad_a[1] ;
    input GND_net;
    input clk_1MHz;
    input clk_1MHz_enable_91;
    output \SLO_buf[0] ;
    input \spi_data_out_r_39__N_4419[0] ;
    output spi_data_out_r_39__N_4197;
    input spi_data_out_r_39__N_4490;
    input n29762;
    output \SLO_buf[29] ;
    output \SLO_buf[28] ;
    output \SLO_buf[27] ;
    output \SLO_buf[26] ;
    output \SLO_buf[25] ;
    output \SLO_buf[24] ;
    output \SLO_buf[23] ;
    output \SLO_buf[22] ;
    output \SLO_buf[21] ;
    output \SLO_buf[20] ;
    output \SLO_buf[19] ;
    output \SLO_buf[18] ;
    output \SLO_buf[17] ;
    output \SLO_buf[16] ;
    output \SLO_buf[15] ;
    output \SLO_buf[14] ;
    output \SLO_buf[9] ;
    output \SLO_buf[8] ;
    output \SLO_buf[7] ;
    output \SLO_buf[6] ;
    output \SLO_buf[5] ;
    output \SLO_buf[4] ;
    output \SLO_buf[3] ;
    output \SLO_buf[2] ;
    output \SLO_buf[1] ;
    output n19351;
    input resetn_c;
    output n29217;
    output n29315;
    input \cs_decoded[2] ;
    input n29306;
    output n8796;
    input OW_ID_N_4464;
    input C_5_c_c;
    output OW_ID_N_4462;
    output reset_r;
    input clk_enable_307;
    input n29097;
    output n1;
    output n1_adj_8;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire MA_Temp_N_4274 /* synthesis is_inv_clock=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    wire clk_1MHz_derived_89 /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz_derived_89 */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire MA_Temp /* synthesis is_clock=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(57[5:12])
    wire [51:0]SLO_buf;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire n29228, n24988;
    wire [7:0]Cnt;   // c:/s_links/sources/slot_cards/stepper.v(62[11:14])
    wire [31:0]n153;
    
    wire n24987;
    wire [11:0]Cnt_NSL;   // c:/s_links/sources/slot_cards/stepper.v(61[12:19])
    wire [11:0]n1290;
    wire [51:0]SLO;   // c:/s_links/sources/slot_cards/stepper.v(63[12:15])
    
    wire clk_1MHz_derived_89_enable_46, clk_1MHz_enable_80;
    wire [7:0]n199;
    
    wire clk_1MHz_derived_89_enable_27, n29148, n4, n19425, n19501, 
        n29250, n28696, n29215, n11851, n29170, n13372, n27453, 
        clk_1MHz_enable_342, NSL, clk_1MHz_enable_100, NSL_N_4485, n24986, 
        n24985, n29312, n19455, n24994, n24993, MA_Temp_N_4277, 
        n28695, n28697, n28694, n24992, n24991, n24990, n24989;
    
    FD1P3IX mode__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_30), .CD(n29239), 
            .CK(clk), .Q(mode[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i2.GSR = "DISABLED";
    FD1P3IX mode__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_30), .CD(n29239), 
            .CK(clk), .Q(mode[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i1.GSR = "DISABLED";
    FD1P3IX digital_output_r_481 (.D(\spi_data_r[0] ), .SP(clk_enable_20), 
            .CD(n29239), .CK(clk), .Q(digital_output_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam digital_output_r_481.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i39 (.D(\SLO_buf[13] ), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i39.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i38 (.D(\SLO_buf[12] ), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i38.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i37 (.D(\SLO_buf[11] ), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i37.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i36 (.D(\SLO_buf[10] ), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i36.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i35 (.D(\spi_data_out_r_39__N_4419[35] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i35.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i34 (.D(\spi_data_out_r_39__N_4419[34] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i34.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i33 (.D(\spi_data_out_r_39__N_4419[33] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i33.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_4419[32] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i31 (.D(SLO_buf[45]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i30 (.D(SLO_buf[44]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i29 (.D(SLO_buf[43]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i28 (.D(SLO_buf[42]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i27 (.D(SLO_buf[41]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i26 (.D(SLO_buf[40]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i25 (.D(SLO_buf[39]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i24 (.D(SLO_buf[38]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i23 (.D(SLO_buf[37]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i22 (.D(SLO_buf[36]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i21 (.D(SLO_buf[35]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i20 (.D(SLO_buf[34]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i19 (.D(SLO_buf[33]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i18 (.D(SLO_buf[32]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i17 (.D(SLO_buf[31]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i16 (.D(SLO_buf[30]), .CK(clk), .CD(n29094), 
            .Q(spi_data_out_r_39__N_4157[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_4419[15] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_4419[14] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_4419[13] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_4419[12] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_4419[11] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_4419[10] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_4419[9] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_4419[8] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_4419[7] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_4419[6] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_4419[5] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_4419[4] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_4419[3] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_4419[2] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_4419[1] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_500 (.A(mode[2]), .B(mode[1]), .Z(n29228)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_500.init = 16'hbbbb;
    LUT4 Select_4099_i1_2_lut_3_lut_4_lut (.A(mode[2]), .B(mode[1]), .C(pin_io_out_19), 
         .D(mode[0]), .Z(\quad_b[1] )) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam Select_4099_i1_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 Select_4092_i1_2_lut_3_lut_4_lut (.A(mode[2]), .B(mode[1]), .C(pin_io_out_18), 
         .D(mode[0]), .Z(\quad_a[1] )) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam Select_4092_i1_2_lut_3_lut_4_lut.init = 16'h0040;
    CCU2D add_552_9 (.A0(Cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24988), 
          .S0(n153[7]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_9.INIT0 = 16'h5aaa;
    defparam add_552_9.INIT1 = 16'h0000;
    defparam add_552_9.INJECT1_0 = "NO";
    defparam add_552_9.INJECT1_1 = "NO";
    CCU2D add_552_7 (.A0(Cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24987), 
          .COUT(n24988), .S0(n153[5]), .S1(n153[6]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_7.INIT0 = 16'h5aaa;
    defparam add_552_7.INIT1 = 16'h5aaa;
    defparam add_552_7.INJECT1_0 = "NO";
    defparam add_552_7.INJECT1_1 = "NO";
    FD1P3IX Cnt_NSL__i0 (.D(n1290[0]), .SP(clk_1MHz_enable_91), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i0.GSR = "DISABLED";
    FD1S3AX SLO_buf_i1 (.D(SLO[0]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i1.GSR = "DISABLED";
    FD1P3AX SLO_i0 (.D(pin_io_out_18), .SP(clk_1MHz_derived_89_enable_46), 
            .CK(clk_1MHz_derived_89), .Q(SLO[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i0 (.D(\spi_data_out_r_39__N_4419[0] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4157[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i0.GSR = "DISABLED";
    FD1S3IX i159_483 (.D(spi_data_out_r_39__N_4490), .CK(clk), .CD(n29239), 
            .Q(spi_data_out_r_39__N_4197)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam i159_483.GSR = "DISABLED";
    FD1P3IX mode__i0 (.D(n29762), .SP(clk_enable_30), .CD(n29239), .CK(clk), 
            .Q(mode[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i0.GSR = "DISABLED";
    FD1P3IX Cnt__i0 (.D(n199[0]), .SP(clk_1MHz_enable_80), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i0.GSR = "DISABLED";
    FD1P3IX SLO_i45 (.D(SLO[44]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i45.GSR = "DISABLED";
    FD1P3IX SLO_i44 (.D(SLO[43]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i44.GSR = "DISABLED";
    FD1P3IX SLO_i43 (.D(SLO[42]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i43.GSR = "DISABLED";
    FD1P3IX SLO_i42 (.D(SLO[41]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i42.GSR = "DISABLED";
    FD1P3IX SLO_i41 (.D(SLO[40]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i41.GSR = "DISABLED";
    FD1P3IX SLO_i40 (.D(SLO[39]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i40.GSR = "DISABLED";
    FD1P3IX SLO_i39 (.D(SLO[38]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i39.GSR = "DISABLED";
    FD1P3IX SLO_i38 (.D(SLO[37]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i38.GSR = "DISABLED";
    FD1P3IX SLO_i37 (.D(SLO[36]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i37.GSR = "DISABLED";
    FD1P3IX SLO_i36 (.D(SLO[35]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i36.GSR = "DISABLED";
    FD1P3IX SLO_i35 (.D(SLO[34]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i35.GSR = "DISABLED";
    FD1P3IX SLO_i34 (.D(SLO[33]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i34.GSR = "DISABLED";
    FD1P3IX SLO_i33 (.D(SLO[32]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i33.GSR = "DISABLED";
    FD1P3IX SLO_i32 (.D(SLO[31]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i32.GSR = "DISABLED";
    FD1P3IX SLO_i31 (.D(SLO[30]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i31.GSR = "DISABLED";
    FD1P3IX SLO_i30 (.D(SLO[29]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i30.GSR = "DISABLED";
    FD1P3IX SLO_i29 (.D(SLO[28]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i29.GSR = "DISABLED";
    FD1P3IX SLO_i28 (.D(SLO[27]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i28.GSR = "DISABLED";
    FD1P3IX SLO_i27 (.D(SLO[26]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i27.GSR = "DISABLED";
    FD1P3IX SLO_i26 (.D(SLO[25]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i26.GSR = "DISABLED";
    FD1P3IX SLO_i25 (.D(SLO[24]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i25.GSR = "DISABLED";
    FD1P3IX SLO_i24 (.D(SLO[23]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i24.GSR = "DISABLED";
    FD1P3IX SLO_i23 (.D(SLO[22]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i23.GSR = "DISABLED";
    FD1P3IX SLO_i22 (.D(SLO[21]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i22.GSR = "DISABLED";
    FD1P3IX SLO_i21 (.D(SLO[20]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i21.GSR = "DISABLED";
    FD1P3IX SLO_i20 (.D(SLO[19]), .SP(clk_1MHz_derived_89_enable_27), .CD(n29148), 
            .CK(clk_1MHz_derived_89), .Q(SLO[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i20.GSR = "DISABLED";
    FD1P3AX SLO_i19 (.D(SLO[18]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i19.GSR = "DISABLED";
    FD1P3AX SLO_i18 (.D(SLO[17]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i18.GSR = "DISABLED";
    FD1P3AX SLO_i17 (.D(SLO[16]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i17.GSR = "DISABLED";
    FD1P3AX SLO_i16 (.D(SLO[15]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i16.GSR = "DISABLED";
    FD1P3AX SLO_i15 (.D(SLO[14]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i15.GSR = "DISABLED";
    FD1P3AX SLO_i14 (.D(SLO[13]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i14.GSR = "DISABLED";
    FD1P3AX SLO_i13 (.D(SLO[12]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i13.GSR = "DISABLED";
    FD1P3AX SLO_i12 (.D(SLO[11]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i12.GSR = "DISABLED";
    FD1P3AX SLO_i11 (.D(SLO[10]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i11.GSR = "DISABLED";
    FD1P3AX SLO_i10 (.D(SLO[9]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i10.GSR = "DISABLED";
    FD1P3AX SLO_i9 (.D(SLO[8]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i9.GSR = "DISABLED";
    FD1P3AX SLO_i8 (.D(SLO[7]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i8.GSR = "DISABLED";
    FD1P3AX SLO_i7 (.D(SLO[6]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i7.GSR = "DISABLED";
    FD1P3AX SLO_i6 (.D(SLO[5]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i6.GSR = "DISABLED";
    FD1P3AX SLO_i5 (.D(SLO[4]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i5.GSR = "DISABLED";
    FD1P3AX SLO_i4 (.D(SLO[3]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i4.GSR = "DISABLED";
    FD1P3AX SLO_i3 (.D(SLO[2]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i3.GSR = "DISABLED";
    FD1P3AX SLO_i2 (.D(SLO[1]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i2.GSR = "DISABLED";
    FD1P3AX SLO_i1 (.D(SLO[0]), .SP(clk_1MHz_derived_89_enable_46), .CK(clk_1MHz_derived_89), 
            .Q(SLO[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i1.GSR = "DISABLED";
    FD1S3AX SLO_buf_i46 (.D(SLO[45]), .CK(MA_Temp_N_4274), .Q(SLO_buf[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i46.GSR = "DISABLED";
    FD1S3AX SLO_buf_i45 (.D(SLO[44]), .CK(MA_Temp_N_4274), .Q(SLO_buf[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i45.GSR = "DISABLED";
    FD1S3AX SLO_buf_i44 (.D(SLO[43]), .CK(MA_Temp_N_4274), .Q(SLO_buf[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i44.GSR = "DISABLED";
    FD1S3AX SLO_buf_i43 (.D(SLO[42]), .CK(MA_Temp_N_4274), .Q(SLO_buf[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i43.GSR = "DISABLED";
    FD1S3AX SLO_buf_i42 (.D(SLO[41]), .CK(MA_Temp_N_4274), .Q(SLO_buf[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i42.GSR = "DISABLED";
    FD1S3AX SLO_buf_i41 (.D(SLO[40]), .CK(MA_Temp_N_4274), .Q(SLO_buf[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i41.GSR = "DISABLED";
    FD1S3AX SLO_buf_i40 (.D(SLO[39]), .CK(MA_Temp_N_4274), .Q(SLO_buf[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i40.GSR = "DISABLED";
    FD1S3AX SLO_buf_i39 (.D(SLO[38]), .CK(MA_Temp_N_4274), .Q(SLO_buf[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i39.GSR = "DISABLED";
    FD1S3AX SLO_buf_i38 (.D(SLO[37]), .CK(MA_Temp_N_4274), .Q(SLO_buf[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i38.GSR = "DISABLED";
    FD1S3AX SLO_buf_i37 (.D(SLO[36]), .CK(MA_Temp_N_4274), .Q(SLO_buf[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i37.GSR = "DISABLED";
    FD1S3AX SLO_buf_i36 (.D(SLO[35]), .CK(MA_Temp_N_4274), .Q(SLO_buf[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i36.GSR = "DISABLED";
    FD1S3AX SLO_buf_i35 (.D(SLO[34]), .CK(MA_Temp_N_4274), .Q(SLO_buf[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i35.GSR = "DISABLED";
    FD1S3AX SLO_buf_i34 (.D(SLO[33]), .CK(MA_Temp_N_4274), .Q(SLO_buf[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i34.GSR = "DISABLED";
    FD1S3AX SLO_buf_i33 (.D(SLO[32]), .CK(MA_Temp_N_4274), .Q(SLO_buf[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i33.GSR = "DISABLED";
    FD1S3AX SLO_buf_i32 (.D(SLO[31]), .CK(MA_Temp_N_4274), .Q(SLO_buf[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i32.GSR = "DISABLED";
    FD1S3AX SLO_buf_i31 (.D(SLO[30]), .CK(MA_Temp_N_4274), .Q(SLO_buf[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i31.GSR = "DISABLED";
    FD1S3AX SLO_buf_i30 (.D(SLO[29]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i30.GSR = "DISABLED";
    FD1S3AX SLO_buf_i29 (.D(SLO[28]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i29.GSR = "DISABLED";
    FD1S3AX SLO_buf_i28 (.D(SLO[27]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i28.GSR = "DISABLED";
    FD1S3AX SLO_buf_i27 (.D(SLO[26]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i27.GSR = "DISABLED";
    FD1S3AX SLO_buf_i26 (.D(SLO[25]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i26.GSR = "DISABLED";
    FD1S3AX SLO_buf_i25 (.D(SLO[24]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i25.GSR = "DISABLED";
    FD1S3AX SLO_buf_i24 (.D(SLO[23]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i24.GSR = "DISABLED";
    FD1S3AX SLO_buf_i23 (.D(SLO[22]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i23.GSR = "DISABLED";
    FD1S3AX SLO_buf_i22 (.D(SLO[21]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i22.GSR = "DISABLED";
    FD1S3AX SLO_buf_i21 (.D(SLO[20]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i21.GSR = "DISABLED";
    FD1S3AX SLO_buf_i20 (.D(SLO[19]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i20.GSR = "DISABLED";
    FD1S3AX SLO_buf_i19 (.D(SLO[18]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i19.GSR = "DISABLED";
    FD1S3AX SLO_buf_i18 (.D(SLO[17]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i18.GSR = "DISABLED";
    FD1S3AX SLO_buf_i17 (.D(SLO[16]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i17.GSR = "DISABLED";
    FD1S3AX SLO_buf_i16 (.D(SLO[15]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i16.GSR = "DISABLED";
    FD1S3AX SLO_buf_i15 (.D(SLO[14]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i15.GSR = "DISABLED";
    FD1S3AX SLO_buf_i14 (.D(SLO[13]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i14.GSR = "DISABLED";
    FD1S3AX SLO_buf_i13 (.D(SLO[12]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i13.GSR = "DISABLED";
    FD1S3AX SLO_buf_i12 (.D(SLO[11]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i12.GSR = "DISABLED";
    FD1S3AX SLO_buf_i11 (.D(SLO[10]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i11.GSR = "DISABLED";
    FD1S3AX SLO_buf_i10 (.D(SLO[9]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i10.GSR = "DISABLED";
    FD1S3AX SLO_buf_i9 (.D(SLO[8]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i9.GSR = "DISABLED";
    FD1P3IX Cnt__i7 (.D(n199[7]), .SP(clk_1MHz_enable_80), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i7.GSR = "DISABLED";
    FD1P3IX Cnt__i6 (.D(n199[6]), .SP(clk_1MHz_enable_80), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i6.GSR = "DISABLED";
    FD1P3IX Cnt__i5 (.D(n199[5]), .SP(clk_1MHz_enable_80), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i5.GSR = "DISABLED";
    FD1P3IX Cnt__i4 (.D(n199[4]), .SP(clk_1MHz_enable_80), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i4.GSR = "DISABLED";
    FD1P3IX Cnt__i3 (.D(n199[3]), .SP(clk_1MHz_enable_80), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i3.GSR = "DISABLED";
    FD1P3IX Cnt__i2 (.D(n199[2]), .SP(clk_1MHz_enable_80), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i1 (.D(n199[1]), .SP(clk_1MHz_enable_80), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i1.GSR = "DISABLED";
    FD1S3AX SLO_buf_i8 (.D(SLO[7]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i8.GSR = "DISABLED";
    FD1S3AX SLO_buf_i7 (.D(SLO[6]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i7.GSR = "DISABLED";
    FD1S3AX SLO_buf_i6 (.D(SLO[5]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i6.GSR = "DISABLED";
    FD1S3AX SLO_buf_i5 (.D(SLO[4]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i5.GSR = "DISABLED";
    FD1S3AX SLO_buf_i4 (.D(SLO[3]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i4.GSR = "DISABLED";
    FD1S3AX SLO_buf_i3 (.D(SLO[2]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i3.GSR = "DISABLED";
    FD1S3AX SLO_buf_i2 (.D(SLO[1]), .CK(MA_Temp_N_4274), .Q(\SLO_buf[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i2.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i11 (.D(n1290[11]), .SP(clk_1MHz_enable_91), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i11.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i10 (.D(n1290[10]), .SP(clk_1MHz_enable_91), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i10.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i9 (.D(n1290[9]), .SP(clk_1MHz_enable_91), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i9.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i8 (.D(n1290[8]), .SP(clk_1MHz_enable_91), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i8.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i7 (.D(n1290[7]), .SP(clk_1MHz_enable_91), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i7.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i6 (.D(n1290[6]), .SP(clk_1MHz_enable_91), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i6.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i5 (.D(n1290[5]), .SP(clk_1MHz_enable_91), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i5.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i4 (.D(n1290[4]), .SP(clk_1MHz_enable_91), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i4.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i3 (.D(n1290[3]), .SP(clk_1MHz_enable_91), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i3.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i2 (.D(n1290[2]), .SP(clk_1MHz_enable_91), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i2.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i1 (.D(n1290[1]), .SP(clk_1MHz_enable_91), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i1.GSR = "DISABLED";
    LUT4 i2_4_lut (.A(Cnt_NSL[11]), .B(Cnt_NSL[9]), .C(Cnt_NSL[10]), .D(n4), 
         .Z(n19351)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'ha080;
    LUT4 i1_2_lut (.A(Cnt_NSL[7]), .B(Cnt_NSL[8]), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i13640_2_lut_3_lut (.A(n19425), .B(n19501), .C(n153[0]), .Z(n199[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13640_2_lut_3_lut.init = 16'h7070;
    LUT4 i13767_2_lut_3_lut (.A(n19425), .B(n19501), .C(n153[7]), .Z(n199[7])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13767_2_lut_3_lut.init = 16'h7070;
    LUT4 i13768_2_lut_3_lut (.A(n19425), .B(n19501), .C(n153[6]), .Z(n199[6])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13768_2_lut_3_lut.init = 16'h7070;
    LUT4 i14298_2_lut_rep_522 (.A(Cnt[4]), .B(Cnt[1]), .Z(n29250)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14298_2_lut_rep_522.init = 16'h8888;
    LUT4 n19425_bdd_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(Cnt[5]), .D(MA_Temp), 
         .Z(n28696)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;
    defparam n19425_bdd_3_lut_4_lut.init = 16'hf708;
    LUT4 i13769_2_lut_3_lut (.A(n19425), .B(n19501), .C(n153[5]), .Z(n199[5])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13769_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(n29215), .D(Cnt[5]), 
         .Z(n11851)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff7;
    LUT4 i13770_2_lut_3_lut (.A(n19425), .B(n19501), .C(n153[4]), .Z(n199[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13770_2_lut_3_lut.init = 16'h7070;
    LUT4 i117_4_lut (.A(n29170), .B(n13372), .C(Cnt[4]), .D(Cnt[1]), 
         .Z(clk_1MHz_derived_89_enable_27)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(132[15:49])
    defparam i117_4_lut.init = 16'h3332;
    LUT4 i13771_2_lut_3_lut (.A(n19425), .B(n19501), .C(n153[3]), .Z(n199[3])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13771_2_lut_3_lut.init = 16'h7070;
    LUT4 i13774_2_lut_3_lut (.A(n19425), .B(n19501), .C(n153[2]), .Z(n199[2])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13774_2_lut_3_lut.init = 16'h7070;
    LUT4 i13775_2_lut_3_lut (.A(n19425), .B(n19501), .C(n153[1]), .Z(n199[1])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13775_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_adj_369 (.A(Cnt[2]), .B(Cnt[3]), .Z(n27453)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_adj_369.init = 16'heeee;
    LUT4 i22848_2_lut_rep_440 (.A(n19351), .B(resetn_c), .Z(clk_1MHz_enable_80)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i22848_2_lut_rep_440.init = 16'hbbbb;
    LUT4 i22616_2_lut_2_lut_3_lut_4_lut (.A(n19351), .B(resetn_c), .C(n19501), 
         .D(n19425), .Z(clk_1MHz_enable_342)) /* synthesis lut_function=(!(A (C (D))+!A (B+(C (D))))) */ ;
    defparam i22616_2_lut_2_lut_3_lut_4_lut.init = 16'h0bbb;
    FD1P3AX NSL_476 (.D(NSL_N_4485), .SP(clk_1MHz_enable_100), .CK(clk_1MHz), 
            .Q(NSL)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam NSL_476.GSR = "DISABLED";
    CCU2D add_552_5 (.A0(Cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24986), 
          .COUT(n24987), .S0(n153[3]), .S1(n153[4]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_5.INIT0 = 16'h5aaa;
    defparam add_552_5.INIT1 = 16'h5aaa;
    defparam add_552_5.INJECT1_0 = "NO";
    defparam add_552_5.INJECT1_1 = "NO";
    CCU2D add_552_3 (.A0(Cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24985), 
          .COUT(n24986), .S0(n153[1]), .S1(n153[2]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_3.INIT0 = 16'h5aaa;
    defparam add_552_3.INIT1 = 16'h5aaa;
    defparam add_552_3.INJECT1_0 = "NO";
    defparam add_552_3.INJECT1_1 = "NO";
    CCU2D add_552_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n24985), 
          .S1(n153[0]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_1.INIT0 = 16'hF000;
    defparam add_552_1.INIT1 = 16'h5555;
    defparam add_552_1.INJECT1_0 = "NO";
    defparam add_552_1.INJECT1_1 = "NO";
    LUT4 i2_4_lut_adj_370 (.A(n29312), .B(Cnt[5]), .C(n13372), .D(n19455), 
         .Z(n19425)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i2_4_lut_adj_370.init = 16'hfefa;
    LUT4 i3_4_lut (.A(n19455), .B(Cnt[5]), .C(n29217), .D(n29312), .Z(n19501)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i14515_4_lut (.A(Cnt[0]), .B(Cnt[4]), .C(n27453), .D(Cnt[1]), 
         .Z(n19455)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i14515_4_lut.init = 16'hc8c0;
    CCU2D add_551_13 (.A0(Cnt_NSL[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n24994), 
          .S0(n1290[11]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_13.INIT0 = 16'h5aaa;
    defparam add_551_13.INIT1 = 16'h0000;
    defparam add_551_13.INJECT1_0 = "NO";
    defparam add_551_13.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_442_4_lut (.A(n27453), .B(Cnt[0]), .C(n29312), .D(Cnt[5]), 
         .Z(n29170)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_rep_442_4_lut.init = 16'hfffe;
    LUT4 Select_4014_i7_3_lut_3_lut_4_lut (.A(mode[0]), .B(n29315), .C(\cs_decoded[2] ), 
         .D(n29306), .Z(n8796)) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam Select_4014_i7_3_lut_3_lut_4_lut.init = 16'hf222;
    CCU2D add_551_11 (.A0(Cnt_NSL[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24993), .COUT(n24994), .S0(n1290[9]), .S1(n1290[10]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_11.INIT0 = 16'h5aaa;
    defparam add_551_11.INIT1 = 16'h5aaa;
    defparam add_551_11.INJECT1_0 = "NO";
    defparam add_551_11.INJECT1_1 = "NO";
    FD1P3IX MA_Temp_474 (.D(MA_Temp_N_4277), .SP(clk_1MHz_enable_342), .CD(n29239), 
            .CK(clk_1MHz), .Q(MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam MA_Temp_474.GSR = "DISABLED";
    LUT4 OW_ID_N_4461_I_0_4_lut (.A(mode[0]), .B(OW_ID_N_4464), .C(n29228), 
         .D(C_5_c_c), .Z(OW_ID_N_4462)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A ((D)+!B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(93[16] 94[93])
    defparam OW_ID_N_4461_I_0_4_lut.init = 16'h0ace;
    FD1P3IX reset_r_480 (.D(n29097), .SP(clk_enable_307), .CD(n29239), 
            .CK(clk), .Q(reset_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam reset_r_480.GSR = "DISABLED";
    PFUMX i23029 (.BLUT(n28696), .ALUT(n28695), .C0(n19501), .Z(n28697));
    LUT4 n28697_bdd_3_lut (.A(n28697), .B(n28694), .C(n29215), .Z(MA_Temp_N_4277)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28697_bdd_3_lut.init = 16'hcaca;
    CCU2D add_551_9 (.A0(Cnt_NSL[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24992), .COUT(n24993), .S0(n1290[7]), .S1(n1290[8]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_9.INIT0 = 16'h5aaa;
    defparam add_551_9.INIT1 = 16'h5aaa;
    defparam add_551_9.INJECT1_0 = "NO";
    defparam add_551_9.INJECT1_1 = "NO";
    CCU2D add_551_7 (.A0(Cnt_NSL[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24991), .COUT(n24992), .S0(n1290[5]), .S1(n1290[6]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_7.INIT0 = 16'h5aaa;
    defparam add_551_7.INIT1 = 16'h5aaa;
    defparam add_551_7.INJECT1_0 = "NO";
    defparam add_551_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_584 (.A(Cnt[7]), .B(Cnt[6]), .Z(n29312)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_rep_584.init = 16'heeee;
    LUT4 i2_3_lut_rep_487_4_lut (.A(Cnt[7]), .B(Cnt[6]), .C(Cnt[0]), .D(n27453), 
         .Z(n29215)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i2_3_lut_rep_487_4_lut.init = 16'hfffe;
    LUT4 n19425_bdd_3_lut_23028 (.A(n19425), .B(n19501), .C(MA_Temp), 
         .Z(n28694)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam n19425_bdd_3_lut_23028.init = 16'h7070;
    LUT4 i1_2_lut_rep_587 (.A(mode[1]), .B(mode[2]), .Z(n29315)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_rep_587.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_489_3_lut (.A(mode[1]), .B(mode[2]), .C(mode[0]), 
         .Z(n29217)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_rep_489_3_lut.init = 16'hbfbf;
    LUT4 n19425_bdd_4_lut_23273 (.A(n19425), .B(n29250), .C(MA_Temp), 
         .D(Cnt[5]), .Z(n28695)) /* synthesis lut_function=(!(A+(B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam n19425_bdd_4_lut_23273.init = 16'h1450;
    LUT4 i1_2_lut_3_lut (.A(mode[1]), .B(mode[2]), .C(mode[0]), .Z(n13372)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_3_lut.init = 16'hfbfb;
    LUT4 Select_3994_i1_2_lut_2_lut_3_lut_4_lut (.A(mode[1]), .B(mode[2]), 
         .C(NSL), .D(mode[0]), .Z(n1)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam Select_3994_i1_2_lut_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 equal_103_i6_1_lut_rep_420_2_lut_3_lut (.A(mode[1]), .B(mode[2]), 
         .C(mode[0]), .Z(n29148)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam equal_103_i6_1_lut_rep_420_2_lut_3_lut.init = 16'h4040;
    LUT4 i4725_2_lut_3_lut_4_lut (.A(mode[1]), .B(mode[2]), .C(clk_1MHz_derived_89_enable_27), 
         .D(mode[0]), .Z(clk_1MHz_derived_89_enable_46)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i4725_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i22628_2_lut_rep_588 (.A(MA_Temp), .B(clk_1MHz), .Z(clk_1MHz_derived_89)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[13:34])
    defparam i22628_2_lut_rep_588.init = 16'h7777;
    LUT4 Select_3991_i1_2_lut_3_lut (.A(MA_Temp), .B(clk_1MHz), .C(mode[2]), 
         .Z(n1_adj_8)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[13:34])
    defparam Select_3991_i1_2_lut_3_lut.init = 16'h7070;
    CCU2D add_551_5 (.A0(Cnt_NSL[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24990), .COUT(n24991), .S0(n1290[3]), .S1(n1290[4]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_5.INIT0 = 16'h5aaa;
    defparam add_551_5.INIT1 = 16'h5aaa;
    defparam add_551_5.INJECT1_0 = "NO";
    defparam add_551_5.INJECT1_1 = "NO";
    CCU2D add_551_3 (.A0(Cnt_NSL[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n24989), .COUT(n24990), .S0(n1290[1]), .S1(n1290[2]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_3.INIT0 = 16'h5aaa;
    defparam add_551_3.INIT1 = 16'h5aaa;
    defparam add_551_3.INJECT1_0 = "NO";
    defparam add_551_3.INJECT1_1 = "NO";
    CCU2D add_551_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n24989), .S1(n1290[0]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_1.INIT0 = 16'hF000;
    defparam add_551_1.INIT1 = 16'h5555;
    defparam add_551_1.INJECT1_0 = "NO";
    defparam add_551_1.INJECT1_1 = "NO";
    LUT4 i14366_3_lut (.A(n19501), .B(resetn_c), .C(n19351), .Z(clk_1MHz_enable_100)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B))) */ ;
    defparam i14366_3_lut.init = 16'h4c4c;
    LUT4 i22625_4_lut (.A(NSL), .B(n19351), .C(n19501), .D(n11851), 
         .Z(NSL_N_4485)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C+(D))))) */ ;
    defparam i22625_4_lut.init = 16'h3b37;
    INV i23374 (.A(MA_Temp), .Z(MA_Temp_N_4274));
    
endmodule
//
// Verilog Description of module \stepper(DEV_ID=5,UART_ADDRESS_WIDTH=4) 
//

module \stepper(DEV_ID=5,UART_ADDRESS_WIDTH=4)  (\SLO_buf[29] , \SLO_buf[28] , 
            \SLO_buf[27] , \SLO_buf[26] , \SLO_buf[25] , \SLO_buf[24] , 
            \SLO_buf[23] , \SLO_buf[22] , \SLO_buf[21] , \SLO_buf[20] , 
            \SLO_buf[19] , \SLO_buf[18] , \SLO_buf[17] , \SLO_buf[16] , 
            \SLO_buf[15] , \SLO_buf[14] , \SLO_buf[13] , \SLO_buf[12] , 
            \SLO_buf[11] , \SLO_buf[10] , \SLO_buf[9] , \SLO_buf[8] , 
            \SLO_buf[7] , \SLO_buf[6] , \SLO_buf[5] , \SLO_buf[4] , 
            \SLO_buf[3] , \SLO_buf[2] , \SLO_buf[1] , clk_1MHz, clk_1MHz_enable_40, 
            n29239, \SLO_buf[0] , pin_io_out_58, spi_data_out_r_39__N_5513, 
            clk, \spi_data_out_r_39__N_5775[0] , mode_adj_7, clk_enable_400, 
            n29762, n19391, spi_data_out_r_39__N_5553, n29108, digital_output_r, 
            clk_enable_199, \spi_data_r[0] , resetn_c, n29301, n29299, 
            \cs_decoded[10] , n8680, n29210, n1, n1_adj_6, reset_r, 
            clk_enable_342, n29075, n29305, \spi_data_out_r_39__N_5775[1] , 
            \spi_data_out_r_39__N_5775[2] , \spi_data_out_r_39__N_5775[3] , 
            \spi_data_out_r_39__N_5775[4] , \spi_data_out_r_39__N_5775[5] , 
            \spi_data_out_r_39__N_5775[6] , \spi_data_out_r_39__N_5775[7] , 
            \spi_data_out_r_39__N_5775[8] , \spi_data_out_r_39__N_5775[9] , 
            \spi_data_out_r_39__N_5775[10] , \spi_data_out_r_39__N_5775[11] , 
            \spi_data_out_r_39__N_5775[12] , \spi_data_out_r_39__N_5775[13] , 
            \spi_data_out_r_39__N_5775[14] , \spi_data_out_r_39__N_5775[15] , 
            \spi_data_out_r_39__N_5775[32] , \spi_data_out_r_39__N_5775[33] , 
            \spi_data_out_r_39__N_5775[34] , \spi_data_out_r_39__N_5775[35] , 
            pin_io_out_59, \quad_b[5] , \quad_a[5] , \spi_data_r[1] , 
            \spi_data_r[2] , mode, n6, n29115, n18550, \spi_addr[1] , 
            \spi_cmd[0] , GND_net) /* synthesis syn_module_defined=1 */ ;
    output \SLO_buf[29] ;
    output \SLO_buf[28] ;
    output \SLO_buf[27] ;
    output \SLO_buf[26] ;
    output \SLO_buf[25] ;
    output \SLO_buf[24] ;
    output \SLO_buf[23] ;
    output \SLO_buf[22] ;
    output \SLO_buf[21] ;
    output \SLO_buf[20] ;
    output \SLO_buf[19] ;
    output \SLO_buf[18] ;
    output \SLO_buf[17] ;
    output \SLO_buf[16] ;
    output \SLO_buf[15] ;
    output \SLO_buf[14] ;
    output \SLO_buf[13] ;
    output \SLO_buf[12] ;
    output \SLO_buf[11] ;
    output \SLO_buf[10] ;
    output \SLO_buf[9] ;
    output \SLO_buf[8] ;
    output \SLO_buf[7] ;
    output \SLO_buf[6] ;
    output \SLO_buf[5] ;
    output \SLO_buf[4] ;
    output \SLO_buf[3] ;
    output \SLO_buf[2] ;
    output \SLO_buf[1] ;
    input clk_1MHz;
    input clk_1MHz_enable_40;
    input n29239;
    output \SLO_buf[0] ;
    input pin_io_out_58;
    output [39:0]spi_data_out_r_39__N_5513;
    input clk;
    input \spi_data_out_r_39__N_5775[0] ;
    output [2:0]mode_adj_7;
    input clk_enable_400;
    input n29762;
    output n19391;
    output spi_data_out_r_39__N_5553;
    input n29108;
    output digital_output_r;
    input clk_enable_199;
    input \spi_data_r[0] ;
    input resetn_c;
    output n29301;
    input n29299;
    input \cs_decoded[10] ;
    output n8680;
    output n29210;
    output n1;
    output n1_adj_6;
    output reset_r;
    input clk_enable_342;
    input n29075;
    output n29305;
    input \spi_data_out_r_39__N_5775[1] ;
    input \spi_data_out_r_39__N_5775[2] ;
    input \spi_data_out_r_39__N_5775[3] ;
    input \spi_data_out_r_39__N_5775[4] ;
    input \spi_data_out_r_39__N_5775[5] ;
    input \spi_data_out_r_39__N_5775[6] ;
    input \spi_data_out_r_39__N_5775[7] ;
    input \spi_data_out_r_39__N_5775[8] ;
    input \spi_data_out_r_39__N_5775[9] ;
    input \spi_data_out_r_39__N_5775[10] ;
    input \spi_data_out_r_39__N_5775[11] ;
    input \spi_data_out_r_39__N_5775[12] ;
    input \spi_data_out_r_39__N_5775[13] ;
    input \spi_data_out_r_39__N_5775[14] ;
    input \spi_data_out_r_39__N_5775[15] ;
    input \spi_data_out_r_39__N_5775[32] ;
    input \spi_data_out_r_39__N_5775[33] ;
    input \spi_data_out_r_39__N_5775[34] ;
    input \spi_data_out_r_39__N_5775[35] ;
    input pin_io_out_59;
    output \quad_b[5] ;
    output \quad_a[5] ;
    input \spi_data_r[1] ;
    input \spi_data_r[2] ;
    input mode;
    output n6;
    input n29115;
    input n18550;
    input \spi_addr[1] ;
    input \spi_cmd[0] ;
    input GND_net;
    
    wire clk_1MHz_derived_277 /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz_derived_277 */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire MA_Temp_N_5630 /* synthesis is_inv_clock=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    wire MA_Temp /* synthesis is_clock=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(57[5:12])
    wire [51:0]SLO;   // c:/s_links/sources/slot_cards/stepper.v(63[12:15])
    
    wire clk_1MHz_derived_277_enable_20, n28867, n28866, n19535, n28868;
    wire [51:0]SLO_buf;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    wire [11:0]Cnt_NSL;   // c:/s_links/sources/slot_cards/stepper.v(61[12:19])
    wire [11:0]n1290;
    wire [7:0]Cnt;   // c:/s_links/sources/slot_cards/stepper.v(62[11:14])
    
    wire clk_1MHz_enable_356;
    wire [7:0]n199;
    
    wire n29166, n13390, clk_1MHz_derived_277_enable_46, n19437;
    wire [31:0]n153;
    
    wire n4, n27456, clk_1MHz_enable_375, clk_1MHz_enable_215, n29280, 
        n29208, n11798, NSL, NSL_N_5841, n29298, MA_Temp_N_5644, 
        n19463, n29088, n28865, MA_Temp_N_5633, n25034, n25033, 
        n25032, n25031, n25030, n25029, n25028, n25027, n25026, 
        n25025;
    
    FD1P3AX SLO_i19 (.D(SLO[18]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i19.GSR = "DISABLED";
    FD1P3AX SLO_i18 (.D(SLO[17]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i18.GSR = "DISABLED";
    FD1P3AX SLO_i17 (.D(SLO[16]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i17.GSR = "DISABLED";
    FD1P3AX SLO_i16 (.D(SLO[15]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i16.GSR = "DISABLED";
    FD1P3AX SLO_i15 (.D(SLO[14]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i15.GSR = "DISABLED";
    FD1P3AX SLO_i14 (.D(SLO[13]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i14.GSR = "DISABLED";
    FD1P3AX SLO_i13 (.D(SLO[12]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i13.GSR = "DISABLED";
    FD1P3AX SLO_i12 (.D(SLO[11]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i12.GSR = "DISABLED";
    FD1P3AX SLO_i11 (.D(SLO[10]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i11.GSR = "DISABLED";
    FD1P3AX SLO_i10 (.D(SLO[9]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i10.GSR = "DISABLED";
    FD1P3AX SLO_i9 (.D(SLO[8]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i9.GSR = "DISABLED";
    FD1P3AX SLO_i8 (.D(SLO[7]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i8.GSR = "DISABLED";
    FD1P3AX SLO_i7 (.D(SLO[6]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i7.GSR = "DISABLED";
    FD1P3AX SLO_i6 (.D(SLO[5]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i6.GSR = "DISABLED";
    FD1P3AX SLO_i5 (.D(SLO[4]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i5.GSR = "DISABLED";
    FD1P3AX SLO_i4 (.D(SLO[3]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i4.GSR = "DISABLED";
    PFUMX i23100 (.BLUT(n28867), .ALUT(n28866), .C0(n19535), .Z(n28868));
    FD1P3AX SLO_i3 (.D(SLO[2]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i3.GSR = "DISABLED";
    FD1P3AX SLO_i2 (.D(SLO[1]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i2.GSR = "DISABLED";
    FD1P3AX SLO_i1 (.D(SLO[0]), .SP(clk_1MHz_derived_277_enable_20), .CK(clk_1MHz_derived_277), 
            .Q(SLO[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i1.GSR = "DISABLED";
    FD1S3AX SLO_buf_i46 (.D(SLO[45]), .CK(MA_Temp_N_5630), .Q(SLO_buf[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i46.GSR = "DISABLED";
    FD1S3AX SLO_buf_i45 (.D(SLO[44]), .CK(MA_Temp_N_5630), .Q(SLO_buf[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i45.GSR = "DISABLED";
    FD1S3AX SLO_buf_i44 (.D(SLO[43]), .CK(MA_Temp_N_5630), .Q(SLO_buf[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i44.GSR = "DISABLED";
    FD1S3AX SLO_buf_i43 (.D(SLO[42]), .CK(MA_Temp_N_5630), .Q(SLO_buf[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i43.GSR = "DISABLED";
    FD1S3AX SLO_buf_i42 (.D(SLO[41]), .CK(MA_Temp_N_5630), .Q(SLO_buf[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i42.GSR = "DISABLED";
    FD1S3AX SLO_buf_i41 (.D(SLO[40]), .CK(MA_Temp_N_5630), .Q(SLO_buf[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i41.GSR = "DISABLED";
    FD1S3AX SLO_buf_i40 (.D(SLO[39]), .CK(MA_Temp_N_5630), .Q(SLO_buf[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i40.GSR = "DISABLED";
    FD1S3AX SLO_buf_i39 (.D(SLO[38]), .CK(MA_Temp_N_5630), .Q(SLO_buf[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i39.GSR = "DISABLED";
    FD1S3AX SLO_buf_i38 (.D(SLO[37]), .CK(MA_Temp_N_5630), .Q(SLO_buf[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i38.GSR = "DISABLED";
    FD1S3AX SLO_buf_i37 (.D(SLO[36]), .CK(MA_Temp_N_5630), .Q(SLO_buf[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i37.GSR = "DISABLED";
    FD1S3AX SLO_buf_i36 (.D(SLO[35]), .CK(MA_Temp_N_5630), .Q(SLO_buf[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i36.GSR = "DISABLED";
    FD1S3AX SLO_buf_i35 (.D(SLO[34]), .CK(MA_Temp_N_5630), .Q(SLO_buf[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i35.GSR = "DISABLED";
    FD1S3AX SLO_buf_i34 (.D(SLO[33]), .CK(MA_Temp_N_5630), .Q(SLO_buf[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i34.GSR = "DISABLED";
    FD1S3AX SLO_buf_i33 (.D(SLO[32]), .CK(MA_Temp_N_5630), .Q(SLO_buf[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i33.GSR = "DISABLED";
    FD1S3AX SLO_buf_i32 (.D(SLO[31]), .CK(MA_Temp_N_5630), .Q(SLO_buf[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i32.GSR = "DISABLED";
    FD1S3AX SLO_buf_i31 (.D(SLO[30]), .CK(MA_Temp_N_5630), .Q(SLO_buf[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i31.GSR = "DISABLED";
    FD1S3AX SLO_buf_i30 (.D(SLO[29]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i30.GSR = "DISABLED";
    FD1S3AX SLO_buf_i29 (.D(SLO[28]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i29.GSR = "DISABLED";
    FD1S3AX SLO_buf_i28 (.D(SLO[27]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i28.GSR = "DISABLED";
    FD1S3AX SLO_buf_i27 (.D(SLO[26]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i27.GSR = "DISABLED";
    FD1S3AX SLO_buf_i26 (.D(SLO[25]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i26.GSR = "DISABLED";
    FD1S3AX SLO_buf_i25 (.D(SLO[24]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i25.GSR = "DISABLED";
    FD1S3AX SLO_buf_i24 (.D(SLO[23]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i24.GSR = "DISABLED";
    FD1S3AX SLO_buf_i23 (.D(SLO[22]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i23.GSR = "DISABLED";
    FD1S3AX SLO_buf_i22 (.D(SLO[21]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i22.GSR = "DISABLED";
    FD1S3AX SLO_buf_i21 (.D(SLO[20]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i21.GSR = "DISABLED";
    FD1S3AX SLO_buf_i20 (.D(SLO[19]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i20.GSR = "DISABLED";
    FD1S3AX SLO_buf_i19 (.D(SLO[18]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i19.GSR = "DISABLED";
    FD1S3AX SLO_buf_i18 (.D(SLO[17]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i18.GSR = "DISABLED";
    FD1S3AX SLO_buf_i17 (.D(SLO[16]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i17.GSR = "DISABLED";
    FD1S3AX SLO_buf_i16 (.D(SLO[15]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i16.GSR = "DISABLED";
    FD1S3AX SLO_buf_i15 (.D(SLO[14]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i15.GSR = "DISABLED";
    FD1S3AX SLO_buf_i14 (.D(SLO[13]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i14.GSR = "DISABLED";
    FD1S3AX SLO_buf_i13 (.D(SLO[12]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i13.GSR = "DISABLED";
    FD1S3AX SLO_buf_i12 (.D(SLO[11]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i12.GSR = "DISABLED";
    FD1S3AX SLO_buf_i11 (.D(SLO[10]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i11.GSR = "DISABLED";
    FD1S3AX SLO_buf_i10 (.D(SLO[9]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i10.GSR = "DISABLED";
    FD1S3AX SLO_buf_i9 (.D(SLO[8]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i9.GSR = "DISABLED";
    FD1S3AX SLO_buf_i8 (.D(SLO[7]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i8.GSR = "DISABLED";
    FD1S3AX SLO_buf_i7 (.D(SLO[6]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i7.GSR = "DISABLED";
    FD1S3AX SLO_buf_i6 (.D(SLO[5]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i6.GSR = "DISABLED";
    FD1S3AX SLO_buf_i5 (.D(SLO[4]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i5.GSR = "DISABLED";
    FD1S3AX SLO_buf_i4 (.D(SLO[3]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i4.GSR = "DISABLED";
    FD1S3AX SLO_buf_i3 (.D(SLO[2]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i3.GSR = "DISABLED";
    FD1S3AX SLO_buf_i2 (.D(SLO[1]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i2.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i11 (.D(n1290[11]), .SP(clk_1MHz_enable_40), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i11.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i10 (.D(n1290[10]), .SP(clk_1MHz_enable_40), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i10.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i9 (.D(n1290[9]), .SP(clk_1MHz_enable_40), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i9.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i8 (.D(n1290[8]), .SP(clk_1MHz_enable_40), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i8.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i7 (.D(n1290[7]), .SP(clk_1MHz_enable_40), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i7.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i6 (.D(n1290[6]), .SP(clk_1MHz_enable_40), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i6.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i5 (.D(n1290[5]), .SP(clk_1MHz_enable_40), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i5.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i4 (.D(n1290[4]), .SP(clk_1MHz_enable_40), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i4.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i3 (.D(n1290[3]), .SP(clk_1MHz_enable_40), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i3.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i2 (.D(n1290[2]), .SP(clk_1MHz_enable_40), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i2.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i1 (.D(n1290[1]), .SP(clk_1MHz_enable_40), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i1.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i0 (.D(n1290[0]), .SP(clk_1MHz_enable_40), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i0.GSR = "DISABLED";
    FD1S3AX SLO_buf_i1 (.D(SLO[0]), .CK(MA_Temp_N_5630), .Q(\SLO_buf[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i1.GSR = "DISABLED";
    FD1P3AX SLO_i0 (.D(pin_io_out_58), .SP(clk_1MHz_derived_277_enable_20), 
            .CK(clk_1MHz_derived_277), .Q(SLO[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i0 (.D(\spi_data_out_r_39__N_5775[0] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i0.GSR = "DISABLED";
    FD1P3IX mode__i0 (.D(n29762), .SP(clk_enable_400), .CD(n29239), .CK(clk), 
            .Q(mode_adj_7[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i0.GSR = "DISABLED";
    FD1P3IX Cnt__i0 (.D(n199[0]), .SP(clk_1MHz_enable_356), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i0.GSR = "DISABLED";
    LUT4 i117_4_lut (.A(n29166), .B(n13390), .C(Cnt[1]), .D(Cnt[4]), 
         .Z(clk_1MHz_derived_277_enable_46)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(132[15:49])
    defparam i117_4_lut.init = 16'h3332;
    LUT4 i13671_2_lut_3_lut (.A(n19437), .B(n19535), .C(n153[0]), .Z(n199[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13671_2_lut_3_lut.init = 16'h7070;
    LUT4 i13699_2_lut_3_lut (.A(n19437), .B(n19535), .C(n153[1]), .Z(n199[1])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13699_2_lut_3_lut.init = 16'h7070;
    LUT4 i13698_2_lut_3_lut (.A(n19437), .B(n19535), .C(n153[2]), .Z(n199[2])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13698_2_lut_3_lut.init = 16'h7070;
    LUT4 i13697_2_lut_3_lut (.A(n19437), .B(n19535), .C(n153[3]), .Z(n199[3])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13697_2_lut_3_lut.init = 16'h7070;
    LUT4 i13696_2_lut_3_lut (.A(n19437), .B(n19535), .C(n153[4]), .Z(n199[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13696_2_lut_3_lut.init = 16'h7070;
    LUT4 i13695_2_lut_3_lut (.A(n19437), .B(n19535), .C(n153[5]), .Z(n199[5])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13695_2_lut_3_lut.init = 16'h7070;
    LUT4 i13694_2_lut_3_lut (.A(n19437), .B(n19535), .C(n153[6]), .Z(n199[6])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13694_2_lut_3_lut.init = 16'h7070;
    LUT4 i13693_2_lut_3_lut (.A(n19437), .B(n19535), .C(n153[7]), .Z(n199[7])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13693_2_lut_3_lut.init = 16'h7070;
    LUT4 i2_4_lut (.A(Cnt_NSL[11]), .B(Cnt_NSL[9]), .C(Cnt_NSL[10]), .D(n4), 
         .Z(n19391)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut.init = 16'ha080;
    LUT4 i1_2_lut (.A(Cnt_NSL[7]), .B(Cnt_NSL[8]), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1S3IX i159_483 (.D(n29108), .CK(clk), .CD(n29239), .Q(spi_data_out_r_39__N_5553)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam i159_483.GSR = "DISABLED";
    LUT4 i1_2_lut_adj_367 (.A(Cnt[2]), .B(Cnt[3]), .Z(n27456)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_adj_367.init = 16'heeee;
    FD1P3IX digital_output_r_481 (.D(\spi_data_r[0] ), .SP(clk_enable_199), 
            .CD(n29239), .CK(clk), .Q(digital_output_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam digital_output_r_481.GSR = "DISABLED";
    LUT4 i22688_2_lut_rep_419 (.A(n19391), .B(resetn_c), .Z(clk_1MHz_enable_356)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i22688_2_lut_rep_419.init = 16'hbbbb;
    LUT4 i22959_2_lut_2_lut_3_lut_4_lut (.A(n19391), .B(resetn_c), .C(n19535), 
         .D(n19437), .Z(clk_1MHz_enable_375)) /* synthesis lut_function=(!(A (C (D))+!A (B+(C (D))))) */ ;
    defparam i22959_2_lut_2_lut_3_lut_4_lut.init = 16'h0bbb;
    LUT4 i14352_3_lut (.A(n19535), .B(resetn_c), .C(n19391), .Z(clk_1MHz_enable_215)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B))) */ ;
    defparam i14352_3_lut.init = 16'h4c4c;
    LUT4 i22883_2_lut_rep_552 (.A(Cnt[4]), .B(Cnt[1]), .Z(n29280)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i22883_2_lut_rep_552.init = 16'h7777;
    LUT4 i1_2_lut_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(n29208), .D(Cnt[5]), 
         .Z(n11798)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff7;
    LUT4 i22662_4_lut (.A(NSL), .B(n19391), .C(n19535), .D(n11798), 
         .Z(NSL_N_5841)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C+(D))))) */ ;
    defparam i22662_4_lut.init = 16'h3b37;
    LUT4 n19437_bdd_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(Cnt[5]), .D(MA_Temp), 
         .Z(n28867)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;
    defparam n19437_bdd_3_lut_4_lut.init = 16'hf708;
    LUT4 i1_2_lut_rep_438_4_lut (.A(n27456), .B(Cnt[0]), .C(n29298), .D(Cnt[5]), 
         .Z(n29166)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_rep_438_4_lut.init = 16'hfffe;
    LUT4 Select_3898_i7_3_lut_4_lut (.A(mode_adj_7[0]), .B(n29301), .C(n29299), 
         .D(\cs_decoded[10] ), .Z(n8680)) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam Select_3898_i7_3_lut_4_lut.init = 16'hf222;
    FD1P3AX NSL_476 (.D(NSL_N_5841), .SP(clk_1MHz_enable_215), .CK(clk_1MHz), 
            .Q(NSL)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam NSL_476.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_570 (.A(Cnt[6]), .B(Cnt[7]), .Z(n29298)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_570.init = 16'heeee;
    LUT4 i2_3_lut_rep_480_4_lut (.A(Cnt[6]), .B(Cnt[7]), .C(Cnt[0]), .D(n27456), 
         .Z(n29208)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_480_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_573 (.A(mode_adj_7[1]), .B(mode_adj_7[2]), .Z(n29301)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_rep_573.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_482_3_lut (.A(mode_adj_7[1]), .B(mode_adj_7[2]), .C(mode_adj_7[0]), 
         .Z(n29210)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_rep_482_3_lut.init = 16'hbfbf;
    LUT4 i4812_2_lut_3_lut_4_lut (.A(mode_adj_7[1]), .B(mode_adj_7[2]), 
         .C(clk_1MHz_derived_277_enable_46), .D(mode_adj_7[0]), .Z(clk_1MHz_derived_277_enable_20)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i4812_2_lut_3_lut_4_lut.init = 16'hf4f0;
    LUT4 i1_2_lut_3_lut (.A(mode_adj_7[1]), .B(mode_adj_7[2]), .C(mode_adj_7[0]), 
         .Z(n13390)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_3_lut.init = 16'hfbfb;
    LUT4 Select_3878_i1_2_lut_3_lut_4_lut (.A(mode_adj_7[1]), .B(mode_adj_7[2]), 
         .C(NSL), .D(mode_adj_7[0]), .Z(n1)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam Select_3878_i1_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 equal_151_i6_1_lut_2_lut_3_lut (.A(mode_adj_7[1]), .B(mode_adj_7[2]), 
         .C(mode_adj_7[0]), .Z(MA_Temp_N_5644)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam equal_151_i6_1_lut_2_lut_3_lut.init = 16'h4040;
    LUT4 i22665_2_lut_rep_574 (.A(MA_Temp), .B(clk_1MHz), .Z(clk_1MHz_derived_277)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[13:34])
    defparam i22665_2_lut_rep_574.init = 16'h7777;
    LUT4 Select_3875_i1_2_lut_3_lut (.A(MA_Temp), .B(clk_1MHz), .C(mode_adj_7[2]), 
         .Z(n1_adj_6)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[13:34])
    defparam Select_3875_i1_2_lut_3_lut.init = 16'h7070;
    LUT4 i2_4_lut_adj_368 (.A(n29298), .B(Cnt[5]), .C(n13390), .D(n19463), 
         .Z(n19437)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i2_4_lut_adj_368.init = 16'hfefa;
    LUT4 i3_4_lut (.A(n19463), .B(Cnt[5]), .C(n29210), .D(n29298), .Z(n19535)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 i14523_4_lut (.A(Cnt[0]), .B(Cnt[4]), .C(n27456), .D(Cnt[1]), 
         .Z(n19463)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i14523_4_lut.init = 16'hc8c0;
    FD1P3IX SLO_i20 (.D(SLO[19]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i20.GSR = "DISABLED";
    FD1P3IX reset_r_480 (.D(n29075), .SP(clk_enable_342), .CD(n29239), 
            .CK(clk), .Q(reset_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam reset_r_480.GSR = "DISABLED";
    FD1P3IX SLO_i21 (.D(SLO[20]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i21.GSR = "DISABLED";
    FD1P3IX SLO_i22 (.D(SLO[21]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i22.GSR = "DISABLED";
    FD1P3IX SLO_i23 (.D(SLO[22]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i23.GSR = "DISABLED";
    FD1P3IX SLO_i24 (.D(SLO[23]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i24.GSR = "DISABLED";
    FD1P3IX SLO_i25 (.D(SLO[24]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i25.GSR = "DISABLED";
    FD1P3IX SLO_i26 (.D(SLO[25]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i26.GSR = "DISABLED";
    FD1P3IX SLO_i27 (.D(SLO[26]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i27.GSR = "DISABLED";
    FD1P3IX SLO_i28 (.D(SLO[27]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i28.GSR = "DISABLED";
    FD1P3IX SLO_i29 (.D(SLO[28]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i29.GSR = "DISABLED";
    FD1P3IX SLO_i30 (.D(SLO[29]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i30.GSR = "DISABLED";
    FD1P3IX SLO_i31 (.D(SLO[30]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i31.GSR = "DISABLED";
    FD1P3IX SLO_i32 (.D(SLO[31]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i32.GSR = "DISABLED";
    FD1P3IX SLO_i33 (.D(SLO[32]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i33.GSR = "DISABLED";
    FD1P3IX SLO_i34 (.D(SLO[33]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i34.GSR = "DISABLED";
    FD1P3IX SLO_i35 (.D(SLO[34]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i35.GSR = "DISABLED";
    FD1P3IX SLO_i36 (.D(SLO[35]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i36.GSR = "DISABLED";
    FD1P3IX SLO_i37 (.D(SLO[36]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i37.GSR = "DISABLED";
    FD1P3IX SLO_i38 (.D(SLO[37]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i38.GSR = "DISABLED";
    FD1P3IX SLO_i39 (.D(SLO[38]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i39.GSR = "DISABLED";
    FD1P3IX SLO_i40 (.D(SLO[39]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i40.GSR = "DISABLED";
    FD1P3IX SLO_i41 (.D(SLO[40]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i41.GSR = "DISABLED";
    FD1P3IX SLO_i42 (.D(SLO[41]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i42.GSR = "DISABLED";
    FD1P3IX SLO_i43 (.D(SLO[42]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i43.GSR = "DISABLED";
    FD1P3IX SLO_i44 (.D(SLO[43]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i44.GSR = "DISABLED";
    FD1P3IX SLO_i45 (.D(SLO[44]), .SP(clk_1MHz_derived_277_enable_46), .CD(MA_Temp_N_5644), 
            .CK(clk_1MHz_derived_277), .Q(SLO[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i45.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_577 (.A(mode_adj_7[0]), .B(mode_adj_7[2]), .Z(n29305)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_577.init = 16'heeee;
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_5775[1] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_5775[2] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_5775[3] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_5775[4] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_5775[5] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_5775[6] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_5775[7] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_5775[8] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_5775[9] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_5775[10] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_5775[11] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_5775[12] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_5775[13] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_5775[14] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_5775[15] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i16 (.D(SLO_buf[30]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i17 (.D(SLO_buf[31]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i18 (.D(SLO_buf[32]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i19 (.D(SLO_buf[33]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i20 (.D(SLO_buf[34]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i21 (.D(SLO_buf[35]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i22 (.D(SLO_buf[36]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i23 (.D(SLO_buf[37]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i24 (.D(SLO_buf[38]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i25 (.D(SLO_buf[39]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i26 (.D(SLO_buf[40]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i27 (.D(SLO_buf[41]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i28 (.D(SLO_buf[42]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i29 (.D(SLO_buf[43]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i30 (.D(SLO_buf[44]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i31 (.D(SLO_buf[45]), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_5775[32] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i33 (.D(\spi_data_out_r_39__N_5775[33] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i33.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i34 (.D(\spi_data_out_r_39__N_5775[34] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i34.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i35 (.D(\spi_data_out_r_39__N_5775[35] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_5513[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i35.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i36 (.D(\SLO_buf[10] ), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i36.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i37 (.D(\SLO_buf[11] ), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i37.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i38 (.D(\SLO_buf[12] ), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i38.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i39 (.D(\SLO_buf[13] ), .CK(clk), .CD(n29088), 
            .Q(spi_data_out_r_39__N_5513[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i39.GSR = "DISABLED";
    LUT4 Select_4095_i1_2_lut_3_lut_4_lut (.A(mode_adj_7[0]), .B(mode_adj_7[2]), 
         .C(pin_io_out_59), .D(mode_adj_7[1]), .Z(\quad_b[5] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam Select_4095_i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 Select_4088_i1_2_lut_3_lut_4_lut (.A(mode_adj_7[0]), .B(mode_adj_7[2]), 
         .C(pin_io_out_58), .D(mode_adj_7[1]), .Z(\quad_a[5] )) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam Select_4088_i1_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 n19437_bdd_3_lut_23099 (.A(n19437), .B(n19535), .C(MA_Temp), 
         .Z(n28865)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam n19437_bdd_3_lut_23099.init = 16'h7070;
    FD1P3IX mode__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_400), .CD(n29239), 
            .CK(clk), .Q(mode_adj_7[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i1.GSR = "DISABLED";
    FD1P3IX mode__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_400), .CD(n29239), 
            .CK(clk), .Q(mode_adj_7[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i1 (.D(n199[1]), .SP(clk_1MHz_enable_356), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i1.GSR = "DISABLED";
    FD1P3IX Cnt__i2 (.D(n199[2]), .SP(clk_1MHz_enable_356), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i3 (.D(n199[3]), .SP(clk_1MHz_enable_356), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i3.GSR = "DISABLED";
    FD1P3IX Cnt__i4 (.D(n199[4]), .SP(clk_1MHz_enable_356), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i4.GSR = "DISABLED";
    FD1P3IX Cnt__i5 (.D(n199[5]), .SP(clk_1MHz_enable_356), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i5.GSR = "DISABLED";
    FD1P3IX Cnt__i6 (.D(n199[6]), .SP(clk_1MHz_enable_356), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i6.GSR = "DISABLED";
    FD1P3IX Cnt__i7 (.D(n199[7]), .SP(clk_1MHz_enable_356), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i7.GSR = "DISABLED";
    LUT4 i2_2_lut_3_lut_4_lut (.A(mode_adj_7[0]), .B(mode_adj_7[2]), .C(mode), 
         .D(mode_adj_7[1]), .Z(n6)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_2_lut_3_lut_4_lut.init = 16'hfffe;
    FD1P3IX MA_Temp_474 (.D(MA_Temp_N_5633), .SP(clk_1MHz_enable_375), .CD(n29239), 
            .CK(clk_1MHz), .Q(MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam MA_Temp_474.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_360_4_lut (.A(n29115), .B(n18550), .C(\spi_addr[1] ), 
         .D(\spi_cmd[0] ), .Z(n29088)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_2_lut_rep_360_4_lut.init = 16'hfffb;
    CCU2D add_551_13 (.A0(Cnt_NSL[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25034), 
          .S0(n1290[11]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_13.INIT0 = 16'h5aaa;
    defparam add_551_13.INIT1 = 16'h0000;
    defparam add_551_13.INJECT1_0 = "NO";
    defparam add_551_13.INJECT1_1 = "NO";
    CCU2D add_551_11 (.A0(Cnt_NSL[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25033), .COUT(n25034), .S0(n1290[9]), .S1(n1290[10]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_11.INIT0 = 16'h5aaa;
    defparam add_551_11.INIT1 = 16'h5aaa;
    defparam add_551_11.INJECT1_0 = "NO";
    defparam add_551_11.INJECT1_1 = "NO";
    CCU2D add_551_9 (.A0(Cnt_NSL[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25032), .COUT(n25033), .S0(n1290[7]), .S1(n1290[8]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_9.INIT0 = 16'h5aaa;
    defparam add_551_9.INIT1 = 16'h5aaa;
    defparam add_551_9.INJECT1_0 = "NO";
    defparam add_551_9.INJECT1_1 = "NO";
    CCU2D add_551_7 (.A0(Cnt_NSL[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25031), .COUT(n25032), .S0(n1290[5]), .S1(n1290[6]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_7.INIT0 = 16'h5aaa;
    defparam add_551_7.INIT1 = 16'h5aaa;
    defparam add_551_7.INJECT1_0 = "NO";
    defparam add_551_7.INJECT1_1 = "NO";
    CCU2D add_551_5 (.A0(Cnt_NSL[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25030), .COUT(n25031), .S0(n1290[3]), .S1(n1290[4]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_5.INIT0 = 16'h5aaa;
    defparam add_551_5.INIT1 = 16'h5aaa;
    defparam add_551_5.INJECT1_0 = "NO";
    defparam add_551_5.INJECT1_1 = "NO";
    CCU2D add_551_3 (.A0(Cnt_NSL[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25029), .COUT(n25030), .S0(n1290[1]), .S1(n1290[2]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_3.INIT0 = 16'h5aaa;
    defparam add_551_3.INIT1 = 16'h5aaa;
    defparam add_551_3.INJECT1_0 = "NO";
    defparam add_551_3.INJECT1_1 = "NO";
    CCU2D add_551_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n25029), .S1(n1290[0]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_1.INIT0 = 16'hF000;
    defparam add_551_1.INIT1 = 16'h5555;
    defparam add_551_1.INJECT1_0 = "NO";
    defparam add_551_1.INJECT1_1 = "NO";
    CCU2D add_552_9 (.A0(Cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25028), 
          .S0(n153[7]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_9.INIT0 = 16'h5aaa;
    defparam add_552_9.INIT1 = 16'h0000;
    defparam add_552_9.INJECT1_0 = "NO";
    defparam add_552_9.INJECT1_1 = "NO";
    CCU2D add_552_7 (.A0(Cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25027), 
          .COUT(n25028), .S0(n153[5]), .S1(n153[6]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_7.INIT0 = 16'h5aaa;
    defparam add_552_7.INIT1 = 16'h5aaa;
    defparam add_552_7.INJECT1_0 = "NO";
    defparam add_552_7.INJECT1_1 = "NO";
    CCU2D add_552_5 (.A0(Cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25026), 
          .COUT(n25027), .S0(n153[3]), .S1(n153[4]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_5.INIT0 = 16'h5aaa;
    defparam add_552_5.INIT1 = 16'h5aaa;
    defparam add_552_5.INJECT1_0 = "NO";
    defparam add_552_5.INJECT1_1 = "NO";
    CCU2D add_552_3 (.A0(Cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25025), 
          .COUT(n25026), .S0(n153[1]), .S1(n153[2]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_3.INIT0 = 16'h5aaa;
    defparam add_552_3.INIT1 = 16'h5aaa;
    defparam add_552_3.INJECT1_0 = "NO";
    defparam add_552_3.INJECT1_1 = "NO";
    CCU2D add_552_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n25025), 
          .S1(n153[0]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_1.INIT0 = 16'hF000;
    defparam add_552_1.INIT1 = 16'h5555;
    defparam add_552_1.INJECT1_0 = "NO";
    defparam add_552_1.INJECT1_1 = "NO";
    LUT4 n19437_bdd_4_lut_23181 (.A(n19437), .B(n29280), .C(MA_Temp), 
         .D(Cnt[5]), .Z(n28866)) /* synthesis lut_function=(!(A+!(B (C)+!B !(C (D)+!C !(D))))) */ ;
    defparam n19437_bdd_4_lut_23181.init = 16'h4150;
    LUT4 n28868_bdd_3_lut (.A(n28868), .B(n28865), .C(n29208), .Z(MA_Temp_N_5633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28868_bdd_3_lut.init = 16'hcaca;
    INV i23369 (.A(MA_Temp), .Z(MA_Temp_N_5630));
    
endmodule
//
// Verilog Description of module \uart_controller(DEV_ID=10,UART_ADDRESS_WIDTH=4) 
//

module \uart_controller(DEV_ID=10,UART_ADDRESS_WIDTH=4)  (C_1_c_0, clk, 
            clk_enable_509, n29239, \spi_data_r[0] , C_2_c_1, \spi_data_r[1] , 
            C_3_c_2, \spi_data_r[2] , C_4_c_3, \spi_data_r[3] ) /* synthesis syn_module_defined=1 */ ;
    output C_1_c_0;
    input clk;
    input clk_enable_509;
    input n29239;
    input \spi_data_r[0] ;
    output C_2_c_1;
    input \spi_data_r[1] ;
    output C_3_c_2;
    input \spi_data_r[2] ;
    output C_4_c_3;
    input \spi_data_r[3] ;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    FD1P3IX uart_slot_en_r__i1 (.D(\spi_data_r[0] ), .SP(clk_enable_509), 
            .CD(n29239), .CK(clk), .Q(C_1_c_0)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=252, LSE_RLINE=263 */ ;   // c:/s_links/sources/uart_controller.v(57[8] 65[4])
    defparam uart_slot_en_r__i1.GSR = "DISABLED";
    FD1P3IX uart_slot_en_r__i2 (.D(\spi_data_r[1] ), .SP(clk_enable_509), 
            .CD(n29239), .CK(clk), .Q(C_2_c_1)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=252, LSE_RLINE=263 */ ;   // c:/s_links/sources/uart_controller.v(57[8] 65[4])
    defparam uart_slot_en_r__i2.GSR = "DISABLED";
    FD1P3IX uart_slot_en_r__i3 (.D(\spi_data_r[2] ), .SP(clk_enable_509), 
            .CD(n29239), .CK(clk), .Q(C_3_c_2)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=252, LSE_RLINE=263 */ ;   // c:/s_links/sources/uart_controller.v(57[8] 65[4])
    defparam uart_slot_en_r__i3.GSR = "DISABLED";
    FD1P3IX uart_slot_en_r__i4 (.D(\spi_data_r[3] ), .SP(clk_enable_509), 
            .CD(n29239), .CK(clk), .Q(C_4_c_3)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=252, LSE_RLINE=263 */ ;   // c:/s_links/sources/uart_controller.v(57[8] 65[4])
    defparam uart_slot_en_r__i4.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \piezo(DEV_ID=5,UART_ADDRESS_WIDTH=4) 
//

module \piezo(DEV_ID=5,UART_ADDRESS_WIDTH=4)  (mode, clk, clk_enable_174, 
            n29239, \spi_data_r[0] , mode_adj_5, digital_output_r, n26523, 
            n29199, mode_adj_3, n6, mode_adj_4, n27186, C_3_c_2, 
            C_4_c_3, n29313, C_2_c_1, C_1_c_0, n29191, \cs_decoded[11] , 
            n2, n8850, C_5_c_c, n26579, n8840) /* synthesis syn_module_defined=1 */ ;
    output mode;
    input clk;
    input clk_enable_174;
    input n29239;
    input \spi_data_r[0] ;
    input [2:0]mode_adj_5;
    input digital_output_r;
    output n26523;
    output n29199;
    input mode_adj_3;
    input n6;
    input mode_adj_4;
    output n27186;
    input C_3_c_2;
    input C_4_c_3;
    output n29313;
    input C_2_c_1;
    input C_1_c_0;
    output n29191;
    input \cs_decoded[11] ;
    output n2;
    output n8850;
    input C_5_c_c;
    output n26579;
    output n8840;
    
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    wire n29263;
    
    FD1P3IX mode_38 (.D(\spi_data_r[0] ), .SP(clk_enable_174), .CD(n29239), 
            .CK(clk), .Q(mode)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=632, LSE_RLINE=661 */ ;   // c:/s_links/sources/slot_cards/piezo.v(55[8] 63[4])
    defparam mode_38.GSR = "DISABLED";
    LUT4 i2_2_lut_rep_535 (.A(mode_adj_5[0]), .B(mode_adj_5[1]), .Z(n29263)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_rep_535.init = 16'h8888;
    LUT4 i3_3_lut_4_lut (.A(mode_adj_5[0]), .B(mode_adj_5[1]), .C(digital_output_r), 
         .D(mode_adj_5[2]), .Z(n26523)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i3_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_4_lut (.A(n29199), .B(mode_adj_3), .C(n6), .D(mode_adj_4), 
         .Z(n27186)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;
    defparam i1_4_lut.init = 16'h5554;
    LUT4 i13790_2_lut_rep_585 (.A(C_3_c_2), .B(C_4_c_3), .Z(n29313)) /* synthesis lut_function=(A (B)) */ ;
    defparam i13790_2_lut_rep_585.init = 16'h8888;
    LUT4 equal_288_i7_2_lut_rep_471_3_lut_4_lut (.A(C_3_c_2), .B(C_4_c_3), 
         .C(C_2_c_1), .D(C_1_c_0), .Z(n29199)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam equal_288_i7_2_lut_rep_471_3_lut_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut_rep_463_3_lut_4_lut (.A(C_3_c_2), .B(C_4_c_3), .C(C_1_c_0), 
         .D(C_2_c_1), .Z(n29191)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_2_lut_rep_463_3_lut_4_lut.init = 16'hff7f;
    LUT4 Select_3891_i2_2_lut (.A(\cs_decoded[11] ), .B(mode), .Z(n2)) /* synthesis lut_function=(A (B)) */ ;
    defparam Select_3891_i2_2_lut.init = 16'h8888;
    LUT4 i4128_1_lut (.A(mode), .Z(n8850)) /* synthesis lut_function=(!(A)) */ ;
    defparam i4128_1_lut.init = 16'h5555;
    LUT4 i22838_4_lut (.A(mode_adj_5[2]), .B(C_5_c_c), .C(n29263), .D(n27186), 
         .Z(n26579)) /* synthesis lut_function=(A (B+!(D))+!A !(B (C)+!B (C+(D)))) */ ;
    defparam i22838_4_lut.init = 16'h8caf;
    LUT4 i1_1_lut (.A(mode_adj_5[2]), .Z(n8840)) /* synthesis lut_function=(!(A)) */ ;
    defparam i1_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module \stepper(DEV_ID=3,UART_ADDRESS_WIDTH=4) 
//

module \stepper(DEV_ID=3,UART_ADDRESS_WIDTH=4)  (mode_adj_2, pin_io_out_38, 
            \quad_a[3] , clk_1MHz, n29239, clk_1MHz_enable_182, n29203, 
            \SLO_buf[0] , spi_data_out_r_39__N_4835, clk, \spi_data_out_r_39__N_5097[0] , 
            clk_enable_86, n29762, \spi_data_r[2] , \spi_data_r[1] , 
            n29093, \SLO_buf[13] , \SLO_buf[12] , \SLO_buf[11] , \SLO_buf[10] , 
            \spi_data_out_r_39__N_5097[35] , \spi_data_out_r_39__N_5097[34] , 
            \spi_data_out_r_39__N_5097[33] , \spi_data_out_r_39__N_5097[32] , 
            \spi_data_out_r_39__N_5097[15] , \spi_data_out_r_39__N_5097[14] , 
            \spi_data_out_r_39__N_5097[13] , \spi_data_out_r_39__N_5097[12] , 
            \spi_data_out_r_39__N_5097[11] , \spi_data_out_r_39__N_5097[10] , 
            \spi_data_out_r_39__N_5097[9] , \spi_data_out_r_39__N_5097[8] , 
            \spi_data_out_r_39__N_5097[7] , \spi_data_out_r_39__N_5097[6] , 
            \spi_data_out_r_39__N_5097[5] , \spi_data_out_r_39__N_5097[4] , 
            \spi_data_out_r_39__N_5097[3] , \spi_data_out_r_39__N_5097[2] , 
            \spi_data_out_r_39__N_5097[1] , n29317, \SLO_buf[29] , \SLO_buf[28] , 
            \SLO_buf[27] , \SLO_buf[26] , \SLO_buf[25] , \SLO_buf[24] , 
            \SLO_buf[23] , \SLO_buf[22] , \SLO_buf[21] , \SLO_buf[20] , 
            \SLO_buf[19] , \SLO_buf[18] , \SLO_buf[17] , \SLO_buf[16] , 
            \SLO_buf[15] , \SLO_buf[14] , \SLO_buf[9] , \SLO_buf[8] , 
            \SLO_buf[7] , \SLO_buf[6] , \SLO_buf[5] , \SLO_buf[4] , 
            \SLO_buf[3] , \SLO_buf[2] , \SLO_buf[1] , digital_output_r, 
            clk_enable_164, \spi_data_r[0] , spi_data_out_r_39__N_4875, 
            n19371, resetn_c, GND_net, NSL, mode, n29300, n29149, 
            pin_io_out_39, \quad_b[3] , reset_r, clk_enable_340, n29110, 
            n1, mode_adj_1, n8716, n29115, \spi_cmd[2] , n13413) /* synthesis syn_module_defined=1 */ ;
    output [2:0]mode_adj_2;
    input pin_io_out_38;
    output \quad_a[3] ;
    input clk_1MHz;
    input n29239;
    input clk_1MHz_enable_182;
    output n29203;
    output \SLO_buf[0] ;
    output [39:0]spi_data_out_r_39__N_4835;
    input clk;
    input \spi_data_out_r_39__N_5097[0] ;
    input clk_enable_86;
    input n29762;
    input \spi_data_r[2] ;
    input \spi_data_r[1] ;
    input n29093;
    output \SLO_buf[13] ;
    output \SLO_buf[12] ;
    output \SLO_buf[11] ;
    output \SLO_buf[10] ;
    input \spi_data_out_r_39__N_5097[35] ;
    input \spi_data_out_r_39__N_5097[34] ;
    input \spi_data_out_r_39__N_5097[33] ;
    input \spi_data_out_r_39__N_5097[32] ;
    input \spi_data_out_r_39__N_5097[15] ;
    input \spi_data_out_r_39__N_5097[14] ;
    input \spi_data_out_r_39__N_5097[13] ;
    input \spi_data_out_r_39__N_5097[12] ;
    input \spi_data_out_r_39__N_5097[11] ;
    input \spi_data_out_r_39__N_5097[10] ;
    input \spi_data_out_r_39__N_5097[9] ;
    input \spi_data_out_r_39__N_5097[8] ;
    input \spi_data_out_r_39__N_5097[7] ;
    input \spi_data_out_r_39__N_5097[6] ;
    input \spi_data_out_r_39__N_5097[5] ;
    input \spi_data_out_r_39__N_5097[4] ;
    input \spi_data_out_r_39__N_5097[3] ;
    input \spi_data_out_r_39__N_5097[2] ;
    input \spi_data_out_r_39__N_5097[1] ;
    output n29317;
    output \SLO_buf[29] ;
    output \SLO_buf[28] ;
    output \SLO_buf[27] ;
    output \SLO_buf[26] ;
    output \SLO_buf[25] ;
    output \SLO_buf[24] ;
    output \SLO_buf[23] ;
    output \SLO_buf[22] ;
    output \SLO_buf[21] ;
    output \SLO_buf[20] ;
    output \SLO_buf[19] ;
    output \SLO_buf[18] ;
    output \SLO_buf[17] ;
    output \SLO_buf[16] ;
    output \SLO_buf[15] ;
    output \SLO_buf[14] ;
    output \SLO_buf[9] ;
    output \SLO_buf[8] ;
    output \SLO_buf[7] ;
    output \SLO_buf[6] ;
    output \SLO_buf[5] ;
    output \SLO_buf[4] ;
    output \SLO_buf[3] ;
    output \SLO_buf[2] ;
    output \SLO_buf[1] ;
    output digital_output_r;
    input clk_enable_164;
    input \spi_data_r[0] ;
    output spi_data_out_r_39__N_4875;
    output n19371;
    input resetn_c;
    input GND_net;
    output NSL;
    input mode;
    input n29300;
    output n29149;
    input pin_io_out_39;
    output \quad_b[3] ;
    output reset_r;
    input clk_enable_340;
    input n29110;
    output n1;
    input mode_adj_1;
    output n8716;
    input n29115;
    input \spi_cmd[2] ;
    input n13413;
    
    wire MA_Temp /* synthesis is_clock=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(57[5:12])
    wire clk_1MHz /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire MA_Temp_N_4952 /* synthesis is_inv_clock=1 */ ;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    wire clk_1MHz_derived_179 /* synthesis is_clock=1, SET_AS_NETWORK=clk_1MHz_derived_179 */ ;   // c:/s_links/sources/mcm_top.v(145[6:14])
    wire clk /* synthesis SET_AS_NETWORK=clk, is_clock=1 */ ;   // c:/s_links/sources/mcm_top.v(79[18:21])
    
    wire clk_1MHz_enable_1, MA_Temp_N_4955;
    wire [11:0]Cnt_NSL;   // c:/s_links/sources/slot_cards/stepper.v(61[12:19])
    wire [11:0]n1290;
    wire [7:0]Cnt;   // c:/s_links/sources/slot_cards/stepper.v(62[11:14])
    
    wire n29223, n28991, n29209, n11824, clk_1MHz_enable_109;
    wire [7:0]n199;
    
    wire n29226, n13369, n29229, n27411;
    wire [51:0]SLO;   // c:/s_links/sources/slot_cards/stepper.v(63[12:15])
    
    wire clk_1MHz_derived_179_enable_46;
    wire [51:0]SLO_buf;   // c:/s_links/sources/slot_cards/stepper.v(64[12:19])
    
    wire clk_1MHz_derived_179_enable_27, n29167, n4, spi_data_out_r_39__N_5168, 
        n19517, n19431, n28992, n28989, n28990, n25014, n25013, 
        clk_1MHz_enable_102, NSL_N_5163, n25012, n25011, n25010, n25009, 
        n25008;
    wire [31:0]n153;
    
    wire n25007, n25006, n25005, n19459;
    
    LUT4 Select_4090_i1_2_lut_4_lut (.A(mode_adj_2[0]), .B(mode_adj_2[1]), 
         .C(mode_adj_2[2]), .D(pin_io_out_38), .Z(\quad_a[3] )) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam Select_4090_i1_2_lut_4_lut.init = 16'h0400;
    FD1P3IX MA_Temp_474 (.D(MA_Temp_N_4955), .SP(clk_1MHz_enable_1), .CD(n29239), 
            .CK(clk_1MHz), .Q(MA_Temp)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam MA_Temp_474.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i0 (.D(n1290[0]), .SP(clk_1MHz_enable_182), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i0.GSR = "DISABLED";
    LUT4 i14324_2_lut_rep_495 (.A(Cnt[4]), .B(Cnt[1]), .Z(n29223)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14324_2_lut_rep_495.init = 16'h8888;
    LUT4 n19431_bdd_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(Cnt[5]), .D(MA_Temp), 
         .Z(n28991)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;
    defparam n19431_bdd_3_lut_4_lut.init = 16'hf708;
    LUT4 i1_2_lut_3_lut_4_lut (.A(Cnt[4]), .B(Cnt[1]), .C(n29209), .D(Cnt[5]), 
         .Z(n11824)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff7;
    FD1P3IX Cnt__i0 (.D(n199[0]), .SP(clk_1MHz_enable_109), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i0.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_498 (.A(mode_adj_2[1]), .B(mode_adj_2[0]), .Z(n29226)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_rep_498.init = 16'heeee;
    LUT4 i1_2_lut_rep_475_3_lut (.A(mode_adj_2[1]), .B(mode_adj_2[0]), .C(mode_adj_2[2]), 
         .Z(n29203)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_rep_475_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut (.A(mode_adj_2[1]), .B(mode_adj_2[0]), .C(mode_adj_2[2]), 
         .Z(n13369)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(111[27:54])
    defparam i1_2_lut_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_501 (.A(Cnt[2]), .B(Cnt[3]), .Z(n29229)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_rep_501.init = 16'heeee;
    LUT4 i2_3_lut_rep_481_4_lut (.A(Cnt[2]), .B(Cnt[3]), .C(n27411), .D(Cnt[0]), 
         .Z(n29209)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i2_3_lut_rep_481_4_lut.init = 16'hfffe;
    FD1S3AX SLO_buf_i1 (.D(SLO[0]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[0] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i1.GSR = "DISABLED";
    FD1P3AX SLO_i0 (.D(pin_io_out_38), .SP(clk_1MHz_derived_179_enable_46), 
            .CK(clk_1MHz_derived_179), .Q(SLO[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i0.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i0 (.D(\spi_data_out_r_39__N_5097[0] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i0.GSR = "DISABLED";
    FD1P3IX mode__i0 (.D(n29762), .SP(clk_enable_86), .CD(n29239), .CK(clk), 
            .Q(mode_adj_2[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i0.GSR = "DISABLED";
    FD1P3IX mode__i2 (.D(\spi_data_r[2] ), .SP(clk_enable_86), .CD(n29239), 
            .CK(clk), .Q(mode_adj_2[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i2.GSR = "DISABLED";
    FD1P3IX mode__i1 (.D(\spi_data_r[1] ), .SP(clk_enable_86), .CD(n29239), 
            .CK(clk), .Q(mode_adj_2[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam mode__i1.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i39 (.D(\SLO_buf[13] ), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i39.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i38 (.D(\SLO_buf[12] ), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i38.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i37 (.D(\SLO_buf[11] ), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i37.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i36 (.D(\SLO_buf[10] ), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i36.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i35 (.D(\spi_data_out_r_39__N_5097[35] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i35.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i34 (.D(\spi_data_out_r_39__N_5097[34] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i34.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i33 (.D(\spi_data_out_r_39__N_5097[33] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i33.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i32 (.D(\spi_data_out_r_39__N_5097[32] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i32.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i31 (.D(SLO_buf[45]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i31.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i30 (.D(SLO_buf[44]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i30.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i29 (.D(SLO_buf[43]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i29.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i28 (.D(SLO_buf[42]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i28.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i27 (.D(SLO_buf[41]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i27.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i26 (.D(SLO_buf[40]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i26.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i25 (.D(SLO_buf[39]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i25.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i24 (.D(SLO_buf[38]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i24.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i23 (.D(SLO_buf[37]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i23.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i22 (.D(SLO_buf[36]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i22.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i21 (.D(SLO_buf[35]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i21.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i20 (.D(SLO_buf[34]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i20.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i19 (.D(SLO_buf[33]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i19.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i18 (.D(SLO_buf[32]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i18.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i17 (.D(SLO_buf[31]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i17.GSR = "DISABLED";
    FD1S3IX spi_data_out_r_i16 (.D(SLO_buf[30]), .CK(clk), .CD(n29093), 
            .Q(spi_data_out_r_39__N_4835[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i16.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i15 (.D(\spi_data_out_r_39__N_5097[15] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i15.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i14 (.D(\spi_data_out_r_39__N_5097[14] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i14.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i13 (.D(\spi_data_out_r_39__N_5097[13] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i13.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i12 (.D(\spi_data_out_r_39__N_5097[12] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i12.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i11 (.D(\spi_data_out_r_39__N_5097[11] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i11.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i10 (.D(\spi_data_out_r_39__N_5097[10] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i10.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i9 (.D(\spi_data_out_r_39__N_5097[9] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i9.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i8 (.D(\spi_data_out_r_39__N_5097[8] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i8.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i7 (.D(\spi_data_out_r_39__N_5097[7] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i7.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i6 (.D(\spi_data_out_r_39__N_5097[6] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i6.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i5 (.D(\spi_data_out_r_39__N_5097[5] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i5.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i4 (.D(\spi_data_out_r_39__N_5097[4] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i4.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i3 (.D(\spi_data_out_r_39__N_5097[3] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i3.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i2 (.D(\spi_data_out_r_39__N_5097[2] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i2.GSR = "DISABLED";
    FD1S3AX spi_data_out_r_i1 (.D(\spi_data_out_r_39__N_5097[1] ), .CK(clk), 
            .Q(spi_data_out_r_39__N_4835[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam spi_data_out_r_i1.GSR = "DISABLED";
    FD1P3IX SLO_i45 (.D(SLO[44]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i45.GSR = "DISABLED";
    FD1P3IX SLO_i44 (.D(SLO[43]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i44.GSR = "DISABLED";
    FD1P3IX SLO_i43 (.D(SLO[42]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i43.GSR = "DISABLED";
    FD1P3IX SLO_i42 (.D(SLO[41]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i42.GSR = "DISABLED";
    FD1P3IX SLO_i41 (.D(SLO[40]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i41.GSR = "DISABLED";
    FD1P3IX SLO_i40 (.D(SLO[39]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i40.GSR = "DISABLED";
    FD1P3IX SLO_i39 (.D(SLO[38]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i39.GSR = "DISABLED";
    FD1P3IX SLO_i38 (.D(SLO[37]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i38.GSR = "DISABLED";
    FD1P3IX SLO_i37 (.D(SLO[36]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i37.GSR = "DISABLED";
    FD1P3IX SLO_i36 (.D(SLO[35]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i36.GSR = "DISABLED";
    FD1P3IX SLO_i35 (.D(SLO[34]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i35.GSR = "DISABLED";
    FD1P3IX SLO_i34 (.D(SLO[33]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i34.GSR = "DISABLED";
    FD1P3IX SLO_i33 (.D(SLO[32]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i33.GSR = "DISABLED";
    FD1P3IX SLO_i32 (.D(SLO[31]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i32.GSR = "DISABLED";
    FD1P3IX SLO_i31 (.D(SLO[30]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i31.GSR = "DISABLED";
    FD1P3IX SLO_i30 (.D(SLO[29]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i30.GSR = "DISABLED";
    FD1P3IX SLO_i29 (.D(SLO[28]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[29])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i29.GSR = "DISABLED";
    FD1P3IX SLO_i28 (.D(SLO[27]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[28])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i28.GSR = "DISABLED";
    FD1P3IX SLO_i27 (.D(SLO[26]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[27])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i27.GSR = "DISABLED";
    FD1P3IX SLO_i26 (.D(SLO[25]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[26])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i26.GSR = "DISABLED";
    FD1P3IX SLO_i25 (.D(SLO[24]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[25])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i25.GSR = "DISABLED";
    FD1P3IX SLO_i24 (.D(SLO[23]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[24])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i24.GSR = "DISABLED";
    FD1P3IX SLO_i23 (.D(SLO[22]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[23])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i23.GSR = "DISABLED";
    FD1P3IX SLO_i22 (.D(SLO[21]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[22])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i22.GSR = "DISABLED";
    FD1P3IX SLO_i21 (.D(SLO[20]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[21])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i21.GSR = "DISABLED";
    FD1P3IX SLO_i20 (.D(SLO[19]), .SP(clk_1MHz_derived_179_enable_27), .CD(n29317), 
            .CK(clk_1MHz_derived_179), .Q(SLO[20])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i20.GSR = "DISABLED";
    FD1P3AX SLO_i19 (.D(SLO[18]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[19])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i19.GSR = "DISABLED";
    FD1P3AX SLO_i18 (.D(SLO[17]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[18])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i18.GSR = "DISABLED";
    FD1P3AX SLO_i17 (.D(SLO[16]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[17])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i17.GSR = "DISABLED";
    FD1P3AX SLO_i16 (.D(SLO[15]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[16])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i16.GSR = "DISABLED";
    FD1P3AX SLO_i15 (.D(SLO[14]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[15])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i15.GSR = "DISABLED";
    FD1P3AX SLO_i14 (.D(SLO[13]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i14.GSR = "DISABLED";
    FD1P3AX SLO_i13 (.D(SLO[12]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i13.GSR = "DISABLED";
    FD1P3AX SLO_i12 (.D(SLO[11]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i12.GSR = "DISABLED";
    FD1P3AX SLO_i11 (.D(SLO[10]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i11.GSR = "DISABLED";
    FD1P3AX SLO_i10 (.D(SLO[9]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i10.GSR = "DISABLED";
    FD1P3AX SLO_i9 (.D(SLO[8]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i9.GSR = "DISABLED";
    FD1P3AX SLO_i8 (.D(SLO[7]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i8.GSR = "DISABLED";
    FD1P3AX SLO_i7 (.D(SLO[6]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i7.GSR = "DISABLED";
    FD1P3AX SLO_i6 (.D(SLO[5]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i6.GSR = "DISABLED";
    FD1P3AX SLO_i5 (.D(SLO[4]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i5.GSR = "DISABLED";
    FD1P3AX SLO_i4 (.D(SLO[3]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i4.GSR = "DISABLED";
    FD1P3AX SLO_i3 (.D(SLO[2]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i3.GSR = "DISABLED";
    FD1P3AX SLO_i2 (.D(SLO[1]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i2.GSR = "DISABLED";
    FD1P3AX SLO_i1 (.D(SLO[0]), .SP(clk_1MHz_derived_179_enable_46), .CK(clk_1MHz_derived_179), 
            .Q(SLO[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(128[8] 135[4])
    defparam SLO_i1.GSR = "DISABLED";
    FD1S3AX SLO_buf_i46 (.D(SLO[45]), .CK(MA_Temp_N_4952), .Q(SLO_buf[45])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i46.GSR = "DISABLED";
    FD1S3AX SLO_buf_i45 (.D(SLO[44]), .CK(MA_Temp_N_4952), .Q(SLO_buf[44])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i45.GSR = "DISABLED";
    FD1S3AX SLO_buf_i44 (.D(SLO[43]), .CK(MA_Temp_N_4952), .Q(SLO_buf[43])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i44.GSR = "DISABLED";
    FD1S3AX SLO_buf_i43 (.D(SLO[42]), .CK(MA_Temp_N_4952), .Q(SLO_buf[42])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i43.GSR = "DISABLED";
    FD1S3AX SLO_buf_i42 (.D(SLO[41]), .CK(MA_Temp_N_4952), .Q(SLO_buf[41])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i42.GSR = "DISABLED";
    FD1S3AX SLO_buf_i41 (.D(SLO[40]), .CK(MA_Temp_N_4952), .Q(SLO_buf[40])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i41.GSR = "DISABLED";
    FD1S3AX SLO_buf_i40 (.D(SLO[39]), .CK(MA_Temp_N_4952), .Q(SLO_buf[39])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i40.GSR = "DISABLED";
    FD1S3AX SLO_buf_i39 (.D(SLO[38]), .CK(MA_Temp_N_4952), .Q(SLO_buf[38])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i39.GSR = "DISABLED";
    FD1S3AX SLO_buf_i38 (.D(SLO[37]), .CK(MA_Temp_N_4952), .Q(SLO_buf[37])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i38.GSR = "DISABLED";
    FD1S3AX SLO_buf_i37 (.D(SLO[36]), .CK(MA_Temp_N_4952), .Q(SLO_buf[36])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i37.GSR = "DISABLED";
    FD1S3AX SLO_buf_i36 (.D(SLO[35]), .CK(MA_Temp_N_4952), .Q(SLO_buf[35])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i36.GSR = "DISABLED";
    FD1S3AX SLO_buf_i35 (.D(SLO[34]), .CK(MA_Temp_N_4952), .Q(SLO_buf[34])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i35.GSR = "DISABLED";
    FD1S3AX SLO_buf_i34 (.D(SLO[33]), .CK(MA_Temp_N_4952), .Q(SLO_buf[33])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i34.GSR = "DISABLED";
    FD1S3AX SLO_buf_i33 (.D(SLO[32]), .CK(MA_Temp_N_4952), .Q(SLO_buf[32])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i33.GSR = "DISABLED";
    FD1S3AX SLO_buf_i32 (.D(SLO[31]), .CK(MA_Temp_N_4952), .Q(SLO_buf[31])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i32.GSR = "DISABLED";
    FD1S3AX SLO_buf_i31 (.D(SLO[30]), .CK(MA_Temp_N_4952), .Q(SLO_buf[30])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i31.GSR = "DISABLED";
    FD1S3AX SLO_buf_i30 (.D(SLO[29]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[29] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i30.GSR = "DISABLED";
    FD1S3AX SLO_buf_i29 (.D(SLO[28]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[28] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i29.GSR = "DISABLED";
    FD1S3AX SLO_buf_i28 (.D(SLO[27]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[27] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i28.GSR = "DISABLED";
    FD1S3AX SLO_buf_i27 (.D(SLO[26]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[26] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i27.GSR = "DISABLED";
    FD1S3AX SLO_buf_i26 (.D(SLO[25]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[25] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i26.GSR = "DISABLED";
    FD1S3AX SLO_buf_i25 (.D(SLO[24]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[24] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i25.GSR = "DISABLED";
    FD1S3AX SLO_buf_i24 (.D(SLO[23]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[23] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i24.GSR = "DISABLED";
    FD1S3AX SLO_buf_i23 (.D(SLO[22]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[22] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i23.GSR = "DISABLED";
    FD1S3AX SLO_buf_i22 (.D(SLO[21]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[21] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i22.GSR = "DISABLED";
    FD1S3AX SLO_buf_i21 (.D(SLO[20]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[20] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i21.GSR = "DISABLED";
    FD1S3AX SLO_buf_i20 (.D(SLO[19]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[19] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i20.GSR = "DISABLED";
    FD1S3AX SLO_buf_i19 (.D(SLO[18]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[18] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i19.GSR = "DISABLED";
    FD1S3AX SLO_buf_i18 (.D(SLO[17]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[17] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i18.GSR = "DISABLED";
    FD1S3AX SLO_buf_i17 (.D(SLO[16]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[16] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i17.GSR = "DISABLED";
    FD1S3AX SLO_buf_i16 (.D(SLO[15]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i16.GSR = "DISABLED";
    FD1S3AX SLO_buf_i15 (.D(SLO[14]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[14] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i15.GSR = "DISABLED";
    FD1S3AX SLO_buf_i14 (.D(SLO[13]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[13] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i14.GSR = "DISABLED";
    FD1S3AX SLO_buf_i13 (.D(SLO[12]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[12] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i13.GSR = "DISABLED";
    FD1S3AX SLO_buf_i12 (.D(SLO[11]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[11] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i12.GSR = "DISABLED";
    FD1S3AX SLO_buf_i11 (.D(SLO[10]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[10] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i11.GSR = "DISABLED";
    FD1S3AX SLO_buf_i10 (.D(SLO[9]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[9] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i10.GSR = "DISABLED";
    FD1S3AX SLO_buf_i9 (.D(SLO[8]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[8] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i9.GSR = "DISABLED";
    FD1S3AX SLO_buf_i8 (.D(SLO[7]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[7] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i8.GSR = "DISABLED";
    FD1S3AX SLO_buf_i7 (.D(SLO[6]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[6] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i7.GSR = "DISABLED";
    FD1S3AX SLO_buf_i6 (.D(SLO[5]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[5] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i6.GSR = "DISABLED";
    FD1S3AX SLO_buf_i5 (.D(SLO[4]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[4] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i5.GSR = "DISABLED";
    FD1S3AX SLO_buf_i4 (.D(SLO[3]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[3] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i4.GSR = "DISABLED";
    FD1S3AX SLO_buf_i3 (.D(SLO[2]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[2] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i3.GSR = "DISABLED";
    FD1S3AX SLO_buf_i2 (.D(SLO[1]), .CK(MA_Temp_N_4952), .Q(\SLO_buf[1] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(124[8] 126[4])
    defparam SLO_buf_i2.GSR = "DISABLED";
    LUT4 i117_4_lut (.A(n29167), .B(n13369), .C(Cnt[1]), .D(Cnt[4]), 
         .Z(clk_1MHz_derived_179_enable_27)) /* synthesis lut_function=(!(A (B)+!A (B+!(C+(D))))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(132[15:49])
    defparam i117_4_lut.init = 16'h3332;
    LUT4 i1_2_lut (.A(Cnt_NSL[7]), .B(Cnt_NSL[8]), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1P3IX digital_output_r_481 (.D(\spi_data_r[0] ), .SP(clk_enable_164), 
            .CD(n29239), .CK(clk), .Q(digital_output_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam digital_output_r_481.GSR = "DISABLED";
    FD1S3IX i159_483 (.D(spi_data_out_r_39__N_5168), .CK(clk), .CD(n29239), 
            .Q(spi_data_out_r_39__N_4875)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(199[8] 209[4])
    defparam i159_483.GSR = "DISABLED";
    LUT4 i22805_2_lut_rep_410 (.A(n19371), .B(resetn_c), .Z(clk_1MHz_enable_109)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i22805_2_lut_rep_410.init = 16'hbbbb;
    LUT4 i22857_2_lut_2_lut_3_lut_4_lut (.A(n19371), .B(resetn_c), .C(n19517), 
         .D(n19431), .Z(clk_1MHz_enable_1)) /* synthesis lut_function=(!(A (C (D))+!A (B+(C (D))))) */ ;
    defparam i22857_2_lut_2_lut_3_lut_4_lut.init = 16'h0bbb;
    LUT4 n28992_bdd_3_lut (.A(n28992), .B(n28989), .C(n29209), .Z(MA_Temp_N_4955)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28992_bdd_3_lut.init = 16'hcaca;
    LUT4 n19431_bdd_4_lut_23352 (.A(n19431), .B(n29223), .C(MA_Temp), 
         .D(Cnt[5]), .Z(n28990)) /* synthesis lut_function=(!(A+(B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam n19431_bdd_4_lut_23352.init = 16'h1450;
    LUT4 n19431_bdd_3_lut_23130 (.A(n19431), .B(n19517), .C(MA_Temp), 
         .Z(n28989)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam n19431_bdd_3_lut_23130.init = 16'h7070;
    CCU2D add_551_13 (.A0(Cnt_NSL[11]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25014), 
          .S0(n1290[11]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_13.INIT0 = 16'h5aaa;
    defparam add_551_13.INIT1 = 16'h0000;
    defparam add_551_13.INJECT1_0 = "NO";
    defparam add_551_13.INJECT1_1 = "NO";
    CCU2D add_551_11 (.A0(Cnt_NSL[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25013), .COUT(n25014), .S0(n1290[9]), .S1(n1290[10]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_11.INIT0 = 16'h5aaa;
    defparam add_551_11.INIT1 = 16'h5aaa;
    defparam add_551_11.INJECT1_0 = "NO";
    defparam add_551_11.INJECT1_1 = "NO";
    FD1P3AX NSL_476 (.D(NSL_N_5163), .SP(clk_1MHz_enable_102), .CK(clk_1MHz), 
            .Q(NSL)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam NSL_476.GSR = "DISABLED";
    FD1P3IX Cnt__i7 (.D(n199[7]), .SP(clk_1MHz_enable_109), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i7.GSR = "DISABLED";
    FD1P3IX Cnt__i6 (.D(n199[6]), .SP(clk_1MHz_enable_109), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i6.GSR = "DISABLED";
    FD1P3IX Cnt__i5 (.D(n199[5]), .SP(clk_1MHz_enable_109), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i5.GSR = "DISABLED";
    FD1P3IX Cnt__i4 (.D(n199[4]), .SP(clk_1MHz_enable_109), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i4.GSR = "DISABLED";
    FD1P3IX Cnt__i3 (.D(n199[3]), .SP(clk_1MHz_enable_109), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i3.GSR = "DISABLED";
    FD1P3IX Cnt__i2 (.D(n199[2]), .SP(clk_1MHz_enable_109), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i2.GSR = "DISABLED";
    FD1P3IX Cnt__i1 (.D(n199[1]), .SP(clk_1MHz_enable_109), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt__i1.GSR = "DISABLED";
    CCU2D add_551_9 (.A0(Cnt_NSL[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25012), .COUT(n25013), .S0(n1290[7]), .S1(n1290[8]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_9.INIT0 = 16'h5aaa;
    defparam add_551_9.INIT1 = 16'h5aaa;
    defparam add_551_9.INJECT1_0 = "NO";
    defparam add_551_9.INJECT1_1 = "NO";
    CCU2D add_551_7 (.A0(Cnt_NSL[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25011), .COUT(n25012), .S0(n1290[5]), .S1(n1290[6]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_7.INIT0 = 16'h5aaa;
    defparam add_551_7.INIT1 = 16'h5aaa;
    defparam add_551_7.INJECT1_0 = "NO";
    defparam add_551_7.INJECT1_1 = "NO";
    CCU2D add_551_5 (.A0(Cnt_NSL[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25010), .COUT(n25011), .S0(n1290[3]), .S1(n1290[4]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_5.INIT0 = 16'h5aaa;
    defparam add_551_5.INIT1 = 16'h5aaa;
    defparam add_551_5.INJECT1_0 = "NO";
    defparam add_551_5.INJECT1_1 = "NO";
    CCU2D add_551_3 (.A0(Cnt_NSL[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n25009), .COUT(n25010), .S0(n1290[1]), .S1(n1290[2]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_3.INIT0 = 16'h5aaa;
    defparam add_551_3.INIT1 = 16'h5aaa;
    defparam add_551_3.INJECT1_0 = "NO";
    defparam add_551_3.INJECT1_1 = "NO";
    CCU2D add_551_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt_NSL[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n25009), .S1(n1290[0]));   // c:/s_links/sources/slot_cards/stepper.v(104[15:26])
    defparam add_551_1.INIT0 = 16'hF000;
    defparam add_551_1.INIT1 = 16'h5555;
    defparam add_551_1.INJECT1_0 = "NO";
    defparam add_551_1.INJECT1_1 = "NO";
    CCU2D add_552_9 (.A0(Cnt[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25008), 
          .S0(n153[7]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_9.INIT0 = 16'h5aaa;
    defparam add_552_9.INIT1 = 16'h0000;
    defparam add_552_9.INJECT1_0 = "NO";
    defparam add_552_9.INJECT1_1 = "NO";
    CCU2D add_552_7 (.A0(Cnt[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25007), 
          .COUT(n25008), .S0(n153[5]), .S1(n153[6]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_7.INIT0 = 16'h5aaa;
    defparam add_552_7.INIT1 = 16'h5aaa;
    defparam add_552_7.INJECT1_0 = "NO";
    defparam add_552_7.INJECT1_1 = "NO";
    CCU2D add_552_5 (.A0(Cnt[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25006), 
          .COUT(n25007), .S0(n153[3]), .S1(n153[4]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_5.INIT0 = 16'h5aaa;
    defparam add_552_5.INIT1 = 16'h5aaa;
    defparam add_552_5.INJECT1_0 = "NO";
    defparam add_552_5.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_421_4_lut (.A(mode_adj_2[2]), .B(n29226), .C(mode), 
         .D(n29300), .Z(n29149)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_rep_421_4_lut.init = 16'hfffe;
    CCU2D add_552_3 (.A0(Cnt[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n25005), 
          .COUT(n25006), .S0(n153[1]), .S1(n153[2]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_3.INIT0 = 16'h5aaa;
    defparam add_552_3.INIT1 = 16'h5aaa;
    defparam add_552_3.INJECT1_0 = "NO";
    defparam add_552_3.INJECT1_1 = "NO";
    CCU2D add_552_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(Cnt[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n25005), 
          .S1(n153[0]));   // c:/s_links/sources/slot_cards/stepper.v(112[11:16])
    defparam add_552_1.INIT0 = 16'hF000;
    defparam add_552_1.INIT1 = 16'h5555;
    defparam add_552_1.INJECT1_0 = "NO";
    defparam add_552_1.INJECT1_1 = "NO";
    FD1P3IX Cnt_NSL__i11 (.D(n1290[11]), .SP(clk_1MHz_enable_182), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i11.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i10 (.D(n1290[10]), .SP(clk_1MHz_enable_182), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i10.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i9 (.D(n1290[9]), .SP(clk_1MHz_enable_182), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i9.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i8 (.D(n1290[8]), .SP(clk_1MHz_enable_182), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i8.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i7 (.D(n1290[7]), .SP(clk_1MHz_enable_182), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i7.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i6 (.D(n1290[6]), .SP(clk_1MHz_enable_182), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i6.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i5 (.D(n1290[5]), .SP(clk_1MHz_enable_182), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i5.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i4 (.D(n1290[4]), .SP(clk_1MHz_enable_182), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i4.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i3 (.D(n1290[3]), .SP(clk_1MHz_enable_182), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i3.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i2 (.D(n1290[2]), .SP(clk_1MHz_enable_182), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i2.GSR = "DISABLED";
    FD1P3IX Cnt_NSL__i1 (.D(n1290[1]), .SP(clk_1MHz_enable_182), .CD(n29239), 
            .CK(clk_1MHz), .Q(Cnt_NSL[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(97[8] 119[4])
    defparam Cnt_NSL__i1.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_439_4_lut (.A(n29229), .B(Cnt[0]), .C(n27411), .D(Cnt[5]), 
         .Z(n29167)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_rep_439_4_lut.init = 16'hfffe;
    LUT4 Select_4097_i1_2_lut_4_lut (.A(mode_adj_2[0]), .B(mode_adj_2[1]), 
         .C(mode_adj_2[2]), .D(pin_io_out_39), .Z(\quad_b[3] )) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam Select_4097_i1_2_lut_4_lut.init = 16'h0400;
    FD1P3IX reset_r_480 (.D(n29110), .SP(clk_enable_340), .CD(n29239), 
            .CK(clk), .Q(reset_r)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=3, LSE_RCOL=2, LSE_LLINE=364, LSE_RLINE=407 */ ;   // c:/s_links/sources/slot_cards/stepper.v(163[8] 195[4])
    defparam reset_r_480.GSR = "DISABLED";
    LUT4 i22647_2_lut_rep_576 (.A(MA_Temp), .B(clk_1MHz), .Z(clk_1MHz_derived_179)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[13:34])
    defparam i22647_2_lut_rep_576.init = 16'h7777;
    LUT4 Select_3932_i1_2_lut_3_lut (.A(MA_Temp), .B(clk_1MHz), .C(mode_adj_2[2]), 
         .Z(n1)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(122[13:34])
    defparam Select_3932_i1_2_lut_3_lut.init = 16'h7070;
    LUT4 i22866_3_lut_rep_589 (.A(mode_adj_2[2]), .B(mode_adj_2[0]), .C(mode_adj_2[1]), 
         .Z(n29317)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(71[15:39])
    defparam i22866_3_lut_rep_589.init = 16'h0808;
    LUT4 i4795_2_lut_4_lut (.A(mode_adj_2[2]), .B(mode_adj_2[0]), .C(mode_adj_2[1]), 
         .D(clk_1MHz_derived_179_enable_27), .Z(clk_1MHz_derived_179_enable_46)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (D)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(71[15:39])
    defparam i4795_2_lut_4_lut.init = 16'hff08;
    LUT4 i22747_2_lut_4_lut (.A(mode_adj_2[2]), .B(mode_adj_2[0]), .C(mode_adj_2[1]), 
         .D(mode_adj_1), .Z(n8716)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(71[15:39])
    defparam i22747_2_lut_4_lut.init = 16'h00f7;
    LUT4 i22650_4_lut (.A(n29093), .B(n29115), .C(\spi_cmd[2] ), .D(n13413), 
         .Z(spi_data_out_r_39__N_5168)) /* synthesis lut_function=(!(A (B+((D)+!C)))) */ ;
    defparam i22650_4_lut.init = 16'h5575;
    LUT4 i2_4_lut (.A(n27411), .B(Cnt[5]), .C(n13369), .D(n19459), .Z(n19431)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i2_4_lut.init = 16'hfefa;
    LUT4 i3_4_lut (.A(n19459), .B(Cnt[5]), .C(n29317), .D(n27411), .Z(n19517)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i3_4_lut.init = 16'hffef;
    LUT4 i1_2_lut_adj_365 (.A(Cnt[6]), .B(Cnt[7]), .Z(n27411)) /* synthesis lut_function=(A+(B)) */ ;   // c:/s_links/sources/slot_cards/stepper.v(113[8:17])
    defparam i1_2_lut_adj_365.init = 16'heeee;
    LUT4 i14519_4_lut (.A(Cnt[0]), .B(Cnt[4]), .C(n29229), .D(Cnt[1]), 
         .Z(n19459)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;
    defparam i14519_4_lut.init = 16'hc8c0;
    LUT4 i13657_2_lut_3_lut (.A(n19431), .B(n19517), .C(n153[0]), .Z(n199[0])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13657_2_lut_3_lut.init = 16'h7070;
    LUT4 i13742_2_lut_3_lut (.A(n19431), .B(n19517), .C(n153[7]), .Z(n199[7])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13742_2_lut_3_lut.init = 16'h7070;
    LUT4 i13743_2_lut_3_lut (.A(n19431), .B(n19517), .C(n153[6]), .Z(n199[6])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13743_2_lut_3_lut.init = 16'h7070;
    LUT4 i13744_2_lut_3_lut (.A(n19431), .B(n19517), .C(n153[5]), .Z(n199[5])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13744_2_lut_3_lut.init = 16'h7070;
    LUT4 i13745_2_lut_3_lut (.A(n19431), .B(n19517), .C(n153[4]), .Z(n199[4])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13745_2_lut_3_lut.init = 16'h7070;
    LUT4 i13746_2_lut_3_lut (.A(n19431), .B(n19517), .C(n153[3]), .Z(n199[3])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13746_2_lut_3_lut.init = 16'h7070;
    LUT4 i13747_2_lut_3_lut (.A(n19431), .B(n19517), .C(n153[2]), .Z(n199[2])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13747_2_lut_3_lut.init = 16'h7070;
    LUT4 i13748_2_lut_3_lut (.A(n19431), .B(n19517), .C(n153[1]), .Z(n199[1])) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13748_2_lut_3_lut.init = 16'h7070;
    LUT4 i2_4_lut_adj_366 (.A(Cnt_NSL[11]), .B(Cnt_NSL[9]), .C(Cnt_NSL[10]), 
         .D(n4), .Z(n19371)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_366.init = 16'ha080;
    LUT4 i14389_3_lut (.A(n19517), .B(resetn_c), .C(n19371), .Z(clk_1MHz_enable_102)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B))) */ ;
    defparam i14389_3_lut.init = 16'h4c4c;
    LUT4 i22644_4_lut (.A(NSL), .B(n19371), .C(n19517), .D(n11824), 
         .Z(NSL_N_5163)) /* synthesis lut_function=(!(A (B (C+!(D)))+!A (B (C+(D))))) */ ;
    defparam i22644_4_lut.init = 16'h3b37;
    PFUMX i23131 (.BLUT(n28991), .ALUT(n28990), .C0(n19517), .Z(n28992));
    INV i23373 (.A(MA_Temp), .Z(MA_Temp_N_4952));
    
endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.12.0.240.2 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.12/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo2c00 -type bram -wp 10 -rp 0011 -data_width 1 -num_rows 2 -rdata_width 1 -read_reg1 outreg -gsr DISABLED -reset_rel async -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr11211211401afe -pmi -lang verilog  */
/* Thu Apr 21 17:03:17 2022 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr11211211401afe (WrAddress, RdAddress, Data, 
    WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [0:0] WrAddress;
    input wire [0:0] RdAddress;
    input wire [0:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [0:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.DATA_WIDTH_B = 1 ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.DATA_WIDTH_A = 1 ;
    DP8KC pmi_ram_dpXbnonesadr11211211401afe_0_0_0 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), 
        .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), 
        .DIA2(scuba_vlo), .DIA1(Data[0]), .DIA0(scuba_vlo), .ADA12(scuba_vlo), 
        .ADA11(scuba_vlo), .ADA10(scuba_vlo), .ADA9(scuba_vlo), .ADA8(scuba_vlo), 
        .ADA7(scuba_vlo), .ADA6(scuba_vlo), .ADA5(scuba_vlo), .ADA4(scuba_vlo), 
        .ADA3(scuba_vlo), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(WrAddress[0]), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo), 
        .ADB12(scuba_vlo), .ADB11(scuba_vlo), .ADB10(scuba_vlo), .ADB9(scuba_vlo), 
        .ADB8(scuba_vlo), .ADB7(scuba_vlo), .ADB6(scuba_vlo), .ADB5(scuba_vlo), 
        .ADB4(scuba_vlo), .ADB3(scuba_vlo), .ADB2(scuba_vlo), .ADB1(scuba_vlo), 
        .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), 
        .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr11211211401afe__PMIP__2__1__1B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr11211211401afe_0_0_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr11211211401afe__PMIP__2__1__1B
    // exemplar attribute pmi_ram_dpXbnonesadr11211211401afe_0_0_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.12.0.240.2 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.12/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo2c00 -type bram -wp 10 -rp 0011 -data_width 91 -num_rows 2048 -rdata_width 91 -read_reg1 outreg -gsr DISABLED -reset_rel async -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr911120489111204811f45a5e -pmi -lang verilog  */
/* Thu Apr 21 17:03:17 2022 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr911120489111204811f45a5e (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [10:0] WrAddress;
    input wire [10:0] RdAddress;
    input wire [90:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [90:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;
    wire raddr10_ff;
    wire mdout1_1_0;
    wire mdout1_0_0;
    wire mdout1_1_1;
    wire mdout1_0_1;
    wire mdout1_1_2;
    wire mdout1_0_2;
    wire mdout1_1_3;
    wire mdout1_0_3;
    wire mdout1_1_4;
    wire mdout1_0_4;
    wire mdout1_1_5;
    wire mdout1_0_5;
    wire mdout1_1_6;
    wire mdout1_0_6;
    wire mdout1_1_7;
    wire mdout1_0_7;
    wire mdout1_1_8;
    wire mdout1_0_8;
    wire mdout1_1_9;
    wire mdout1_0_9;
    wire mdout1_1_10;
    wire mdout1_0_10;
    wire mdout1_1_11;
    wire mdout1_0_11;
    wire mdout1_1_12;
    wire mdout1_0_12;
    wire mdout1_1_13;
    wire mdout1_0_13;
    wire mdout1_1_14;
    wire mdout1_0_14;
    wire mdout1_1_15;
    wire mdout1_0_15;
    wire mdout1_1_16;
    wire mdout1_0_16;
    wire mdout1_1_17;
    wire mdout1_0_17;
    wire mdout1_1_18;
    wire mdout1_0_18;
    wire mdout1_1_19;
    wire mdout1_0_19;
    wire mdout1_1_20;
    wire mdout1_0_20;
    wire mdout1_1_21;
    wire mdout1_0_21;
    wire mdout1_1_22;
    wire mdout1_0_22;
    wire mdout1_1_23;
    wire mdout1_0_23;
    wire mdout1_1_24;
    wire mdout1_0_24;
    wire mdout1_1_25;
    wire mdout1_0_25;
    wire mdout1_1_26;
    wire mdout1_0_26;
    wire mdout1_1_27;
    wire mdout1_0_27;
    wire mdout1_1_28;
    wire mdout1_0_28;
    wire mdout1_1_29;
    wire mdout1_0_29;
    wire mdout1_1_30;
    wire mdout1_0_30;
    wire mdout1_1_31;
    wire mdout1_0_31;
    wire mdout1_1_32;
    wire mdout1_0_32;
    wire mdout1_1_33;
    wire mdout1_0_33;
    wire mdout1_1_34;
    wire mdout1_0_34;
    wire mdout1_1_35;
    wire mdout1_0_35;
    wire mdout1_1_36;
    wire mdout1_0_36;
    wire mdout1_1_37;
    wire mdout1_0_37;
    wire mdout1_1_38;
    wire mdout1_0_38;
    wire mdout1_1_39;
    wire mdout1_0_39;
    wire mdout1_1_40;
    wire mdout1_0_40;
    wire mdout1_1_41;
    wire mdout1_0_41;
    wire mdout1_1_42;
    wire mdout1_0_42;
    wire mdout1_1_43;
    wire mdout1_0_43;
    wire mdout1_1_44;
    wire mdout1_0_44;
    wire mdout1_1_45;
    wire mdout1_0_45;
    wire mdout1_1_46;
    wire mdout1_0_46;
    wire mdout1_1_47;
    wire mdout1_0_47;
    wire mdout1_1_48;
    wire mdout1_0_48;
    wire mdout1_1_49;
    wire mdout1_0_49;
    wire mdout1_1_50;
    wire mdout1_0_50;
    wire mdout1_1_51;
    wire mdout1_0_51;
    wire mdout1_1_52;
    wire mdout1_0_52;
    wire mdout1_1_53;
    wire mdout1_0_53;
    wire mdout1_1_54;
    wire mdout1_0_54;
    wire mdout1_1_55;
    wire mdout1_0_55;
    wire mdout1_1_56;
    wire mdout1_0_56;
    wire mdout1_1_57;
    wire mdout1_0_57;
    wire mdout1_1_58;
    wire mdout1_0_58;
    wire mdout1_1_59;
    wire mdout1_0_59;
    wire mdout1_1_60;
    wire mdout1_0_60;
    wire mdout1_1_61;
    wire mdout1_0_61;
    wire mdout1_1_62;
    wire mdout1_0_62;
    wire mdout1_1_63;
    wire mdout1_0_63;
    wire mdout1_1_64;
    wire mdout1_0_64;
    wire mdout1_1_65;
    wire mdout1_0_65;
    wire mdout1_1_66;
    wire mdout1_0_66;
    wire mdout1_1_67;
    wire mdout1_0_67;
    wire mdout1_1_68;
    wire mdout1_0_68;
    wire mdout1_1_69;
    wire mdout1_0_69;
    wire mdout1_1_70;
    wire mdout1_0_70;
    wire mdout1_1_71;
    wire mdout1_0_71;
    wire mdout1_1_72;
    wire mdout1_0_72;
    wire mdout1_1_73;
    wire mdout1_0_73;
    wire mdout1_1_74;
    wire mdout1_0_74;
    wire mdout1_1_75;
    wire mdout1_0_75;
    wire mdout1_1_76;
    wire mdout1_0_76;
    wire mdout1_1_77;
    wire mdout1_0_77;
    wire mdout1_1_78;
    wire mdout1_0_78;
    wire mdout1_1_79;
    wire mdout1_0_79;
    wire mdout1_1_80;
    wire mdout1_0_80;
    wire mdout1_1_81;
    wire mdout1_0_81;
    wire mdout1_1_82;
    wire mdout1_0_82;
    wire mdout1_1_83;
    wire mdout1_0_83;
    wire mdout1_1_84;
    wire mdout1_0_84;
    wire mdout1_1_85;
    wire mdout1_0_85;
    wire mdout1_1_86;
    wire mdout1_0_86;
    wire mdout1_1_87;
    wire mdout1_0_87;
    wire mdout1_1_88;
    wire mdout1_0_88;
    wire mdout1_1_89;
    wire mdout1_0_89;
    wire raddr10_ff2;
    wire mdout1_1_90;
    wire mdout1_0_90;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_8), .DOB7(mdout1_0_7), .DOB6(mdout1_0_6), 
        .DOB5(mdout1_0_5), .DOB4(mdout1_0_4), .DOB3(mdout1_0_3), .DOB2(mdout1_0_2), 
        .DOB1(mdout1_0_1), .DOB0(mdout1_0_0))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_17), .DOB7(mdout1_0_16), .DOB6(mdout1_0_15), 
        .DOB5(mdout1_0_14), .DOB4(mdout1_0_13), .DOB3(mdout1_0_12), .DOB2(mdout1_0_11), 
        .DOB1(mdout1_0_10), .DOB0(mdout1_0_9))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_26), .DOB7(mdout1_0_25), .DOB6(mdout1_0_24), 
        .DOB5(mdout1_0_23), .DOB4(mdout1_0_22), .DOB3(mdout1_0_21), .DOB2(mdout1_0_20), 
        .DOB1(mdout1_0_19), .DOB0(mdout1_0_18))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_35), .DOB7(mdout1_0_34), .DOB6(mdout1_0_33), 
        .DOB5(mdout1_0_32), .DOB4(mdout1_0_31), .DOB3(mdout1_0_30), .DOB2(mdout1_0_29), 
        .DOB1(mdout1_0_28), .DOB0(mdout1_0_27))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_44), .DOB7(mdout1_0_43), .DOB6(mdout1_0_42), 
        .DOB5(mdout1_0_41), .DOB4(mdout1_0_40), .DOB3(mdout1_0_39), .DOB2(mdout1_0_38), 
        .DOB1(mdout1_0_37), .DOB0(mdout1_0_36))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_53), .DOB7(mdout1_0_52), .DOB6(mdout1_0_51), 
        .DOB5(mdout1_0_50), .DOB4(mdout1_0_49), .DOB3(mdout1_0_48), .DOB2(mdout1_0_47), 
        .DOB1(mdout1_0_46), .DOB0(mdout1_0_45))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_62), .DOB7(mdout1_0_61), .DOB6(mdout1_0_60), 
        .DOB5(mdout1_0_59), .DOB4(mdout1_0_58), .DOB3(mdout1_0_57), .DOB2(mdout1_0_56), 
        .DOB1(mdout1_0_55), .DOB0(mdout1_0_54))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_71), .DOB7(mdout1_0_70), .DOB6(mdout1_0_69), 
        .DOB5(mdout1_0_68), .DOB4(mdout1_0_67), .DOB3(mdout1_0_66), .DOB2(mdout1_0_65), 
        .DOB1(mdout1_0_64), .DOB0(mdout1_0_63))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_80), .DOB7(mdout1_0_79), .DOB6(mdout1_0_78), 
        .DOB5(mdout1_0_77), .DOB4(mdout1_0_76), .DOB3(mdout1_0_75), .DOB2(mdout1_0_74), 
        .DOB1(mdout1_0_73), .DOB0(mdout1_0_72))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_89), .DOB7(mdout1_0_88), .DOB6(mdout1_0_87), 
        .DOB5(mdout1_0_86), .DOB4(mdout1_0_85), .DOB3(mdout1_0_84), .DOB2(mdout1_0_83), 
        .DOB1(mdout1_0_82), .DOB0(mdout1_0_81))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(), .DOB0(mdout1_0_90))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_8), .DOB7(mdout1_1_7), .DOB6(mdout1_1_6), 
        .DOB5(mdout1_1_5), .DOB4(mdout1_1_4), .DOB3(mdout1_1_3), .DOB2(mdout1_1_2), 
        .DOB1(mdout1_1_1), .DOB0(mdout1_1_0))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_17), .DOB7(mdout1_1_16), .DOB6(mdout1_1_15), 
        .DOB5(mdout1_1_14), .DOB4(mdout1_1_13), .DOB3(mdout1_1_12), .DOB2(mdout1_1_11), 
        .DOB1(mdout1_1_10), .DOB0(mdout1_1_9))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_26), .DOB7(mdout1_1_25), .DOB6(mdout1_1_24), 
        .DOB5(mdout1_1_23), .DOB4(mdout1_1_22), .DOB3(mdout1_1_21), .DOB2(mdout1_1_20), 
        .DOB1(mdout1_1_19), .DOB0(mdout1_1_18))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_35), .DOB7(mdout1_1_34), .DOB6(mdout1_1_33), 
        .DOB5(mdout1_1_32), .DOB4(mdout1_1_31), .DOB3(mdout1_1_30), .DOB2(mdout1_1_29), 
        .DOB1(mdout1_1_28), .DOB0(mdout1_1_27))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_44), .DOB7(mdout1_1_43), .DOB6(mdout1_1_42), 
        .DOB5(mdout1_1_41), .DOB4(mdout1_1_40), .DOB3(mdout1_1_39), .DOB2(mdout1_1_38), 
        .DOB1(mdout1_1_37), .DOB0(mdout1_1_36))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_53), .DOB7(mdout1_1_52), .DOB6(mdout1_1_51), 
        .DOB5(mdout1_1_50), .DOB4(mdout1_1_49), .DOB3(mdout1_1_48), .DOB2(mdout1_1_47), 
        .DOB1(mdout1_1_46), .DOB0(mdout1_1_45))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_62), .DOB7(mdout1_1_61), .DOB6(mdout1_1_60), 
        .DOB5(mdout1_1_59), .DOB4(mdout1_1_58), .DOB3(mdout1_1_57), .DOB2(mdout1_1_56), 
        .DOB1(mdout1_1_55), .DOB0(mdout1_1_54))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_71), .DOB7(mdout1_1_70), .DOB6(mdout1_1_69), 
        .DOB5(mdout1_1_68), .DOB4(mdout1_1_67), .DOB3(mdout1_1_66), .DOB2(mdout1_1_65), 
        .DOB1(mdout1_1_64), .DOB0(mdout1_1_63))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_80), .DOB7(mdout1_1_79), .DOB6(mdout1_1_78), 
        .DOB5(mdout1_1_77), .DOB4(mdout1_1_76), .DOB3(mdout1_1_75), .DOB2(mdout1_1_74), 
        .DOB1(mdout1_1_73), .DOB0(mdout1_1_72))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_89), .DOB7(mdout1_1_88), .DOB6(mdout1_1_87), 
        .DOB5(mdout1_1_86), .DOB4(mdout1_1_85), .DOB3(mdout1_1_84), .DOB2(mdout1_1_83), 
        .DOB1(mdout1_1_82), .DOB0(mdout1_1_81))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(), .DOB0(mdout1_1_90))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    FD1P3DX FF_1 (.D(RdAddress[10]), .SP(RdClockEn), .CK(RdClock), .CD(scuba_vlo), 
        .Q(raddr10_ff))
             /* synthesis GSR="ENABLED" */;

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    FD1P3DX FF_0 (.D(raddr10_ff), .SP(RdClockEn), .CK(RdClock), .CD(scuba_vlo), 
        .Q(raddr10_ff2))
             /* synthesis GSR="ENABLED" */;

    MUX21 mux_90 (.D0(mdout1_0_0), .D1(mdout1_1_0), .SD(raddr10_ff2), .Z(Q[0]));

    MUX21 mux_89 (.D0(mdout1_0_1), .D1(mdout1_1_1), .SD(raddr10_ff2), .Z(Q[1]));

    MUX21 mux_88 (.D0(mdout1_0_2), .D1(mdout1_1_2), .SD(raddr10_ff2), .Z(Q[2]));

    MUX21 mux_87 (.D0(mdout1_0_3), .D1(mdout1_1_3), .SD(raddr10_ff2), .Z(Q[3]));

    MUX21 mux_86 (.D0(mdout1_0_4), .D1(mdout1_1_4), .SD(raddr10_ff2), .Z(Q[4]));

    MUX21 mux_85 (.D0(mdout1_0_5), .D1(mdout1_1_5), .SD(raddr10_ff2), .Z(Q[5]));

    MUX21 mux_84 (.D0(mdout1_0_6), .D1(mdout1_1_6), .SD(raddr10_ff2), .Z(Q[6]));

    MUX21 mux_83 (.D0(mdout1_0_7), .D1(mdout1_1_7), .SD(raddr10_ff2), .Z(Q[7]));

    MUX21 mux_82 (.D0(mdout1_0_8), .D1(mdout1_1_8), .SD(raddr10_ff2), .Z(Q[8]));

    MUX21 mux_81 (.D0(mdout1_0_9), .D1(mdout1_1_9), .SD(raddr10_ff2), .Z(Q[9]));

    MUX21 mux_80 (.D0(mdout1_0_10), .D1(mdout1_1_10), .SD(raddr10_ff2), 
        .Z(Q[10]));

    MUX21 mux_79 (.D0(mdout1_0_11), .D1(mdout1_1_11), .SD(raddr10_ff2), 
        .Z(Q[11]));

    MUX21 mux_78 (.D0(mdout1_0_12), .D1(mdout1_1_12), .SD(raddr10_ff2), 
        .Z(Q[12]));

    MUX21 mux_77 (.D0(mdout1_0_13), .D1(mdout1_1_13), .SD(raddr10_ff2), 
        .Z(Q[13]));

    MUX21 mux_76 (.D0(mdout1_0_14), .D1(mdout1_1_14), .SD(raddr10_ff2), 
        .Z(Q[14]));

    MUX21 mux_75 (.D0(mdout1_0_15), .D1(mdout1_1_15), .SD(raddr10_ff2), 
        .Z(Q[15]));

    MUX21 mux_74 (.D0(mdout1_0_16), .D1(mdout1_1_16), .SD(raddr10_ff2), 
        .Z(Q[16]));

    MUX21 mux_73 (.D0(mdout1_0_17), .D1(mdout1_1_17), .SD(raddr10_ff2), 
        .Z(Q[17]));

    MUX21 mux_72 (.D0(mdout1_0_18), .D1(mdout1_1_18), .SD(raddr10_ff2), 
        .Z(Q[18]));

    MUX21 mux_71 (.D0(mdout1_0_19), .D1(mdout1_1_19), .SD(raddr10_ff2), 
        .Z(Q[19]));

    MUX21 mux_70 (.D0(mdout1_0_20), .D1(mdout1_1_20), .SD(raddr10_ff2), 
        .Z(Q[20]));

    MUX21 mux_69 (.D0(mdout1_0_21), .D1(mdout1_1_21), .SD(raddr10_ff2), 
        .Z(Q[21]));

    MUX21 mux_68 (.D0(mdout1_0_22), .D1(mdout1_1_22), .SD(raddr10_ff2), 
        .Z(Q[22]));

    MUX21 mux_67 (.D0(mdout1_0_23), .D1(mdout1_1_23), .SD(raddr10_ff2), 
        .Z(Q[23]));

    MUX21 mux_66 (.D0(mdout1_0_24), .D1(mdout1_1_24), .SD(raddr10_ff2), 
        .Z(Q[24]));

    MUX21 mux_65 (.D0(mdout1_0_25), .D1(mdout1_1_25), .SD(raddr10_ff2), 
        .Z(Q[25]));

    MUX21 mux_64 (.D0(mdout1_0_26), .D1(mdout1_1_26), .SD(raddr10_ff2), 
        .Z(Q[26]));

    MUX21 mux_63 (.D0(mdout1_0_27), .D1(mdout1_1_27), .SD(raddr10_ff2), 
        .Z(Q[27]));

    MUX21 mux_62 (.D0(mdout1_0_28), .D1(mdout1_1_28), .SD(raddr10_ff2), 
        .Z(Q[28]));

    MUX21 mux_61 (.D0(mdout1_0_29), .D1(mdout1_1_29), .SD(raddr10_ff2), 
        .Z(Q[29]));

    MUX21 mux_60 (.D0(mdout1_0_30), .D1(mdout1_1_30), .SD(raddr10_ff2), 
        .Z(Q[30]));

    MUX21 mux_59 (.D0(mdout1_0_31), .D1(mdout1_1_31), .SD(raddr10_ff2), 
        .Z(Q[31]));

    MUX21 mux_58 (.D0(mdout1_0_32), .D1(mdout1_1_32), .SD(raddr10_ff2), 
        .Z(Q[32]));

    MUX21 mux_57 (.D0(mdout1_0_33), .D1(mdout1_1_33), .SD(raddr10_ff2), 
        .Z(Q[33]));

    MUX21 mux_56 (.D0(mdout1_0_34), .D1(mdout1_1_34), .SD(raddr10_ff2), 
        .Z(Q[34]));

    MUX21 mux_55 (.D0(mdout1_0_35), .D1(mdout1_1_35), .SD(raddr10_ff2), 
        .Z(Q[35]));

    MUX21 mux_54 (.D0(mdout1_0_36), .D1(mdout1_1_36), .SD(raddr10_ff2), 
        .Z(Q[36]));

    MUX21 mux_53 (.D0(mdout1_0_37), .D1(mdout1_1_37), .SD(raddr10_ff2), 
        .Z(Q[37]));

    MUX21 mux_52 (.D0(mdout1_0_38), .D1(mdout1_1_38), .SD(raddr10_ff2), 
        .Z(Q[38]));

    MUX21 mux_51 (.D0(mdout1_0_39), .D1(mdout1_1_39), .SD(raddr10_ff2), 
        .Z(Q[39]));

    MUX21 mux_50 (.D0(mdout1_0_40), .D1(mdout1_1_40), .SD(raddr10_ff2), 
        .Z(Q[40]));

    MUX21 mux_49 (.D0(mdout1_0_41), .D1(mdout1_1_41), .SD(raddr10_ff2), 
        .Z(Q[41]));

    MUX21 mux_48 (.D0(mdout1_0_42), .D1(mdout1_1_42), .SD(raddr10_ff2), 
        .Z(Q[42]));

    MUX21 mux_47 (.D0(mdout1_0_43), .D1(mdout1_1_43), .SD(raddr10_ff2), 
        .Z(Q[43]));

    MUX21 mux_46 (.D0(mdout1_0_44), .D1(mdout1_1_44), .SD(raddr10_ff2), 
        .Z(Q[44]));

    MUX21 mux_45 (.D0(mdout1_0_45), .D1(mdout1_1_45), .SD(raddr10_ff2), 
        .Z(Q[45]));

    MUX21 mux_44 (.D0(mdout1_0_46), .D1(mdout1_1_46), .SD(raddr10_ff2), 
        .Z(Q[46]));

    MUX21 mux_43 (.D0(mdout1_0_47), .D1(mdout1_1_47), .SD(raddr10_ff2), 
        .Z(Q[47]));

    MUX21 mux_42 (.D0(mdout1_0_48), .D1(mdout1_1_48), .SD(raddr10_ff2), 
        .Z(Q[48]));

    MUX21 mux_41 (.D0(mdout1_0_49), .D1(mdout1_1_49), .SD(raddr10_ff2), 
        .Z(Q[49]));

    MUX21 mux_40 (.D0(mdout1_0_50), .D1(mdout1_1_50), .SD(raddr10_ff2), 
        .Z(Q[50]));

    MUX21 mux_39 (.D0(mdout1_0_51), .D1(mdout1_1_51), .SD(raddr10_ff2), 
        .Z(Q[51]));

    MUX21 mux_38 (.D0(mdout1_0_52), .D1(mdout1_1_52), .SD(raddr10_ff2), 
        .Z(Q[52]));

    MUX21 mux_37 (.D0(mdout1_0_53), .D1(mdout1_1_53), .SD(raddr10_ff2), 
        .Z(Q[53]));

    MUX21 mux_36 (.D0(mdout1_0_54), .D1(mdout1_1_54), .SD(raddr10_ff2), 
        .Z(Q[54]));

    MUX21 mux_35 (.D0(mdout1_0_55), .D1(mdout1_1_55), .SD(raddr10_ff2), 
        .Z(Q[55]));

    MUX21 mux_34 (.D0(mdout1_0_56), .D1(mdout1_1_56), .SD(raddr10_ff2), 
        .Z(Q[56]));

    MUX21 mux_33 (.D0(mdout1_0_57), .D1(mdout1_1_57), .SD(raddr10_ff2), 
        .Z(Q[57]));

    MUX21 mux_32 (.D0(mdout1_0_58), .D1(mdout1_1_58), .SD(raddr10_ff2), 
        .Z(Q[58]));

    MUX21 mux_31 (.D0(mdout1_0_59), .D1(mdout1_1_59), .SD(raddr10_ff2), 
        .Z(Q[59]));

    MUX21 mux_30 (.D0(mdout1_0_60), .D1(mdout1_1_60), .SD(raddr10_ff2), 
        .Z(Q[60]));

    MUX21 mux_29 (.D0(mdout1_0_61), .D1(mdout1_1_61), .SD(raddr10_ff2), 
        .Z(Q[61]));

    MUX21 mux_28 (.D0(mdout1_0_62), .D1(mdout1_1_62), .SD(raddr10_ff2), 
        .Z(Q[62]));

    MUX21 mux_27 (.D0(mdout1_0_63), .D1(mdout1_1_63), .SD(raddr10_ff2), 
        .Z(Q[63]));

    MUX21 mux_26 (.D0(mdout1_0_64), .D1(mdout1_1_64), .SD(raddr10_ff2), 
        .Z(Q[64]));

    MUX21 mux_25 (.D0(mdout1_0_65), .D1(mdout1_1_65), .SD(raddr10_ff2), 
        .Z(Q[65]));

    MUX21 mux_24 (.D0(mdout1_0_66), .D1(mdout1_1_66), .SD(raddr10_ff2), 
        .Z(Q[66]));

    MUX21 mux_23 (.D0(mdout1_0_67), .D1(mdout1_1_67), .SD(raddr10_ff2), 
        .Z(Q[67]));

    MUX21 mux_22 (.D0(mdout1_0_68), .D1(mdout1_1_68), .SD(raddr10_ff2), 
        .Z(Q[68]));

    MUX21 mux_21 (.D0(mdout1_0_69), .D1(mdout1_1_69), .SD(raddr10_ff2), 
        .Z(Q[69]));

    MUX21 mux_20 (.D0(mdout1_0_70), .D1(mdout1_1_70), .SD(raddr10_ff2), 
        .Z(Q[70]));

    MUX21 mux_19 (.D0(mdout1_0_71), .D1(mdout1_1_71), .SD(raddr10_ff2), 
        .Z(Q[71]));

    MUX21 mux_18 (.D0(mdout1_0_72), .D1(mdout1_1_72), .SD(raddr10_ff2), 
        .Z(Q[72]));

    MUX21 mux_17 (.D0(mdout1_0_73), .D1(mdout1_1_73), .SD(raddr10_ff2), 
        .Z(Q[73]));

    MUX21 mux_16 (.D0(mdout1_0_74), .D1(mdout1_1_74), .SD(raddr10_ff2), 
        .Z(Q[74]));

    MUX21 mux_15 (.D0(mdout1_0_75), .D1(mdout1_1_75), .SD(raddr10_ff2), 
        .Z(Q[75]));

    MUX21 mux_14 (.D0(mdout1_0_76), .D1(mdout1_1_76), .SD(raddr10_ff2), 
        .Z(Q[76]));

    MUX21 mux_13 (.D0(mdout1_0_77), .D1(mdout1_1_77), .SD(raddr10_ff2), 
        .Z(Q[77]));

    MUX21 mux_12 (.D0(mdout1_0_78), .D1(mdout1_1_78), .SD(raddr10_ff2), 
        .Z(Q[78]));

    MUX21 mux_11 (.D0(mdout1_0_79), .D1(mdout1_1_79), .SD(raddr10_ff2), 
        .Z(Q[79]));

    MUX21 mux_10 (.D0(mdout1_0_80), .D1(mdout1_1_80), .SD(raddr10_ff2), 
        .Z(Q[80]));

    MUX21 mux_9 (.D0(mdout1_0_81), .D1(mdout1_1_81), .SD(raddr10_ff2), .Z(Q[81]));

    MUX21 mux_8 (.D0(mdout1_0_82), .D1(mdout1_1_82), .SD(raddr10_ff2), .Z(Q[82]));

    MUX21 mux_7 (.D0(mdout1_0_83), .D1(mdout1_1_83), .SD(raddr10_ff2), .Z(Q[83]));

    MUX21 mux_6 (.D0(mdout1_0_84), .D1(mdout1_1_84), .SD(raddr10_ff2), .Z(Q[84]));

    MUX21 mux_5 (.D0(mdout1_0_85), .D1(mdout1_1_85), .SD(raddr10_ff2), .Z(Q[85]));

    MUX21 mux_4 (.D0(mdout1_0_86), .D1(mdout1_1_86), .SD(raddr10_ff2), .Z(Q[86]));

    MUX21 mux_3 (.D0(mdout1_0_87), .D1(mdout1_1_87), .SD(raddr10_ff2), .Z(Q[87]));

    MUX21 mux_2 (.D0(mdout1_0_88), .D1(mdout1_1_88), .SD(raddr10_ff2), .Z(Q[88]));

    MUX21 mux_1 (.D0(mdout1_0_89), .D1(mdout1_1_89), .SD(raddr10_ff2), .Z(Q[89]));

    MUX21 mux_0 (.D0(mdout1_0_90), .D1(mdout1_1_90), .SD(raddr10_ff2), .Z(Q[90]));



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0 MEM_INIT_FILE 
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.12.0.240.2 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.12/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo2c00 -type bram -wp 10 -rp 0011 -data_width 1 -num_rows 2 -rdata_width 1 -read_reg1 outreg -gsr DISABLED -reset_rel async -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr11211211401afe -pmi -lang verilog  */
/* Fri Apr 22 14:02:28 2022 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr11211211401afe (WrAddress, RdAddress, Data, 
    WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [0:0] WrAddress;
    input wire [0:0] RdAddress;
    input wire [0:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [0:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.DATA_WIDTH_B = 1 ;
    defparam pmi_ram_dpXbnonesadr11211211401afe_0_0_0.DATA_WIDTH_A = 1 ;
    DP8KC pmi_ram_dpXbnonesadr11211211401afe_0_0_0 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), 
        .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), 
        .DIA2(scuba_vlo), .DIA1(Data[0]), .DIA0(scuba_vlo), .ADA12(scuba_vlo), 
        .ADA11(scuba_vlo), .ADA10(scuba_vlo), .ADA9(scuba_vlo), .ADA8(scuba_vlo), 
        .ADA7(scuba_vlo), .ADA6(scuba_vlo), .ADA5(scuba_vlo), .ADA4(scuba_vlo), 
        .ADA3(scuba_vlo), .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(WrAddress[0]), 
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), 
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB8(scuba_vlo), 
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), 
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo), 
        .ADB12(scuba_vlo), .ADB11(scuba_vlo), .ADB10(scuba_vlo), .ADB9(scuba_vlo), 
        .ADB8(scuba_vlo), .ADB7(scuba_vlo), .ADB6(scuba_vlo), .ADB5(scuba_vlo), 
        .ADB4(scuba_vlo), .ADB3(scuba_vlo), .ADB2(scuba_vlo), .ADB1(scuba_vlo), 
        .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), 
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), 
        .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), 
        .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), 
        .DOB3(), .DOB2(), .DOB1(), .DOB0(Q[0]))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr11211211401afe__PMIP__2__1__1B" */
             /* synthesis MEM_INIT_FILE="" */;



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr11211211401afe_0_0_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr11211211401afe__PMIP__2__1__1B
    // exemplar attribute pmi_ram_dpXbnonesadr11211211401afe_0_0_0 MEM_INIT_FILE 
    // exemplar end

endmodule
/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.12.0.240.2 */
/* Module Version: 6.5 */
/* C:/lscc/diamond/3.12/ispfpga/bin/nt64/scuba -w -bus_exp 7 -bb -arch xo2c00 -type bram -wp 10 -rp 0011 -data_width 91 -num_rows 2048 -rdata_width 91 -read_reg1 outreg -gsr DISABLED -reset_rel async -memformat bin -cascade -1 -n pmi_ram_dpXbnonesadr911120489111204811f45a5e -pmi -lang verilog  */
/* Fri Apr 22 14:02:28 2022 */


`timescale 1 ns / 1 ps
module pmi_ram_dpXbnonesadr911120489111204811f45a5e (WrAddress, 
    RdAddress, Data, WE, RdClock, RdClockEn, Reset, WrClock, WrClockEn, 
    Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [10:0] WrAddress;
    input wire [10:0] RdAddress;
    input wire [90:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [90:0] Q;

    wire scuba_vhi;
    wire scuba_vlo;
    wire raddr10_ff;
    wire mdout1_1_0;
    wire mdout1_0_0;
    wire mdout1_1_1;
    wire mdout1_0_1;
    wire mdout1_1_2;
    wire mdout1_0_2;
    wire mdout1_1_3;
    wire mdout1_0_3;
    wire mdout1_1_4;
    wire mdout1_0_4;
    wire mdout1_1_5;
    wire mdout1_0_5;
    wire mdout1_1_6;
    wire mdout1_0_6;
    wire mdout1_1_7;
    wire mdout1_0_7;
    wire mdout1_1_8;
    wire mdout1_0_8;
    wire mdout1_1_9;
    wire mdout1_0_9;
    wire mdout1_1_10;
    wire mdout1_0_10;
    wire mdout1_1_11;
    wire mdout1_0_11;
    wire mdout1_1_12;
    wire mdout1_0_12;
    wire mdout1_1_13;
    wire mdout1_0_13;
    wire mdout1_1_14;
    wire mdout1_0_14;
    wire mdout1_1_15;
    wire mdout1_0_15;
    wire mdout1_1_16;
    wire mdout1_0_16;
    wire mdout1_1_17;
    wire mdout1_0_17;
    wire mdout1_1_18;
    wire mdout1_0_18;
    wire mdout1_1_19;
    wire mdout1_0_19;
    wire mdout1_1_20;
    wire mdout1_0_20;
    wire mdout1_1_21;
    wire mdout1_0_21;
    wire mdout1_1_22;
    wire mdout1_0_22;
    wire mdout1_1_23;
    wire mdout1_0_23;
    wire mdout1_1_24;
    wire mdout1_0_24;
    wire mdout1_1_25;
    wire mdout1_0_25;
    wire mdout1_1_26;
    wire mdout1_0_26;
    wire mdout1_1_27;
    wire mdout1_0_27;
    wire mdout1_1_28;
    wire mdout1_0_28;
    wire mdout1_1_29;
    wire mdout1_0_29;
    wire mdout1_1_30;
    wire mdout1_0_30;
    wire mdout1_1_31;
    wire mdout1_0_31;
    wire mdout1_1_32;
    wire mdout1_0_32;
    wire mdout1_1_33;
    wire mdout1_0_33;
    wire mdout1_1_34;
    wire mdout1_0_34;
    wire mdout1_1_35;
    wire mdout1_0_35;
    wire mdout1_1_36;
    wire mdout1_0_36;
    wire mdout1_1_37;
    wire mdout1_0_37;
    wire mdout1_1_38;
    wire mdout1_0_38;
    wire mdout1_1_39;
    wire mdout1_0_39;
    wire mdout1_1_40;
    wire mdout1_0_40;
    wire mdout1_1_41;
    wire mdout1_0_41;
    wire mdout1_1_42;
    wire mdout1_0_42;
    wire mdout1_1_43;
    wire mdout1_0_43;
    wire mdout1_1_44;
    wire mdout1_0_44;
    wire mdout1_1_45;
    wire mdout1_0_45;
    wire mdout1_1_46;
    wire mdout1_0_46;
    wire mdout1_1_47;
    wire mdout1_0_47;
    wire mdout1_1_48;
    wire mdout1_0_48;
    wire mdout1_1_49;
    wire mdout1_0_49;
    wire mdout1_1_50;
    wire mdout1_0_50;
    wire mdout1_1_51;
    wire mdout1_0_51;
    wire mdout1_1_52;
    wire mdout1_0_52;
    wire mdout1_1_53;
    wire mdout1_0_53;
    wire mdout1_1_54;
    wire mdout1_0_54;
    wire mdout1_1_55;
    wire mdout1_0_55;
    wire mdout1_1_56;
    wire mdout1_0_56;
    wire mdout1_1_57;
    wire mdout1_0_57;
    wire mdout1_1_58;
    wire mdout1_0_58;
    wire mdout1_1_59;
    wire mdout1_0_59;
    wire mdout1_1_60;
    wire mdout1_0_60;
    wire mdout1_1_61;
    wire mdout1_0_61;
    wire mdout1_1_62;
    wire mdout1_0_62;
    wire mdout1_1_63;
    wire mdout1_0_63;
    wire mdout1_1_64;
    wire mdout1_0_64;
    wire mdout1_1_65;
    wire mdout1_0_65;
    wire mdout1_1_66;
    wire mdout1_0_66;
    wire mdout1_1_67;
    wire mdout1_0_67;
    wire mdout1_1_68;
    wire mdout1_0_68;
    wire mdout1_1_69;
    wire mdout1_0_69;
    wire mdout1_1_70;
    wire mdout1_0_70;
    wire mdout1_1_71;
    wire mdout1_0_71;
    wire mdout1_1_72;
    wire mdout1_0_72;
    wire mdout1_1_73;
    wire mdout1_0_73;
    wire mdout1_1_74;
    wire mdout1_0_74;
    wire mdout1_1_75;
    wire mdout1_0_75;
    wire mdout1_1_76;
    wire mdout1_0_76;
    wire mdout1_1_77;
    wire mdout1_0_77;
    wire mdout1_1_78;
    wire mdout1_0_78;
    wire mdout1_1_79;
    wire mdout1_0_79;
    wire mdout1_1_80;
    wire mdout1_0_80;
    wire mdout1_1_81;
    wire mdout1_0_81;
    wire mdout1_1_82;
    wire mdout1_0_82;
    wire mdout1_1_83;
    wire mdout1_0_83;
    wire mdout1_1_84;
    wire mdout1_0_84;
    wire mdout1_1_85;
    wire mdout1_0_85;
    wire mdout1_1_86;
    wire mdout1_0_86;
    wire mdout1_1_87;
    wire mdout1_0_87;
    wire mdout1_1_88;
    wire mdout1_0_88;
    wire mdout1_1_89;
    wire mdout1_0_89;
    wire raddr10_ff2;
    wire mdout1_1_90;
    wire mdout1_0_90;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_8), .DOB7(mdout1_0_7), .DOB6(mdout1_0_6), 
        .DOB5(mdout1_0_5), .DOB4(mdout1_0_4), .DOB3(mdout1_0_3), .DOB2(mdout1_0_2), 
        .DOB1(mdout1_0_1), .DOB0(mdout1_0_0))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_17), .DOB7(mdout1_0_16), .DOB6(mdout1_0_15), 
        .DOB5(mdout1_0_14), .DOB4(mdout1_0_13), .DOB3(mdout1_0_12), .DOB2(mdout1_0_11), 
        .DOB1(mdout1_0_10), .DOB0(mdout1_0_9))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_26), .DOB7(mdout1_0_25), .DOB6(mdout1_0_24), 
        .DOB5(mdout1_0_23), .DOB4(mdout1_0_22), .DOB3(mdout1_0_21), .DOB2(mdout1_0_20), 
        .DOB1(mdout1_0_19), .DOB0(mdout1_0_18))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_35), .DOB7(mdout1_0_34), .DOB6(mdout1_0_33), 
        .DOB5(mdout1_0_32), .DOB4(mdout1_0_31), .DOB3(mdout1_0_30), .DOB2(mdout1_0_29), 
        .DOB1(mdout1_0_28), .DOB0(mdout1_0_27))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_44), .DOB7(mdout1_0_43), .DOB6(mdout1_0_42), 
        .DOB5(mdout1_0_41), .DOB4(mdout1_0_40), .DOB3(mdout1_0_39), .DOB2(mdout1_0_38), 
        .DOB1(mdout1_0_37), .DOB0(mdout1_0_36))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_53), .DOB7(mdout1_0_52), .DOB6(mdout1_0_51), 
        .DOB5(mdout1_0_50), .DOB4(mdout1_0_49), .DOB3(mdout1_0_48), .DOB2(mdout1_0_47), 
        .DOB1(mdout1_0_46), .DOB0(mdout1_0_45))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_62), .DOB7(mdout1_0_61), .DOB6(mdout1_0_60), 
        .DOB5(mdout1_0_59), .DOB4(mdout1_0_58), .DOB3(mdout1_0_57), .DOB2(mdout1_0_56), 
        .DOB1(mdout1_0_55), .DOB0(mdout1_0_54))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_71), .DOB7(mdout1_0_70), .DOB6(mdout1_0_69), 
        .DOB5(mdout1_0_68), .DOB4(mdout1_0_67), .DOB3(mdout1_0_66), .DOB2(mdout1_0_65), 
        .DOB1(mdout1_0_64), .DOB0(mdout1_0_63))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_80), .DOB7(mdout1_0_79), .DOB6(mdout1_0_78), 
        .DOB5(mdout1_0_77), .DOB4(mdout1_0_76), .DOB3(mdout1_0_75), .DOB2(mdout1_0_74), 
        .DOB1(mdout1_0_73), .DOB0(mdout1_0_72))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_0_89), .DOB7(mdout1_0_88), .DOB6(mdout1_0_87), 
        .DOB5(mdout1_0_86), .DOB4(mdout1_0_85), .DOB3(mdout1_0_84), .DOB2(mdout1_0_83), 
        .DOB1(mdout1_0_82), .DOB0(mdout1_0_81))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.CSDECODE_B = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.CSDECODE_A = "0b000" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(), .DOB0(mdout1_0_90))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10 (.DIA8(Data[8]), 
        .DIA7(Data[7]), .DIA6(Data[6]), .DIA5(Data[5]), .DIA4(Data[4]), 
        .DIA3(Data[3]), .DIA2(Data[2]), .DIA1(Data[1]), .DIA0(Data[0]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_8), .DOB7(mdout1_1_7), .DOB6(mdout1_1_6), 
        .DOB5(mdout1_1_5), .DOB4(mdout1_1_4), .DOB3(mdout1_1_3), .DOB2(mdout1_1_2), 
        .DOB1(mdout1_1_1), .DOB0(mdout1_1_0))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9 (.DIA8(Data[17]), 
        .DIA7(Data[16]), .DIA6(Data[15]), .DIA5(Data[14]), .DIA4(Data[13]), 
        .DIA3(Data[12]), .DIA2(Data[11]), .DIA1(Data[10]), .DIA0(Data[9]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_17), .DOB7(mdout1_1_16), .DOB6(mdout1_1_15), 
        .DOB5(mdout1_1_14), .DOB4(mdout1_1_13), .DOB3(mdout1_1_12), .DOB2(mdout1_1_11), 
        .DOB1(mdout1_1_10), .DOB0(mdout1_1_9))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8 (.DIA8(Data[26]), 
        .DIA7(Data[25]), .DIA6(Data[24]), .DIA5(Data[23]), .DIA4(Data[22]), 
        .DIA3(Data[21]), .DIA2(Data[20]), .DIA1(Data[19]), .DIA0(Data[18]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_26), .DOB7(mdout1_1_25), .DOB6(mdout1_1_24), 
        .DOB5(mdout1_1_23), .DOB4(mdout1_1_22), .DOB3(mdout1_1_21), .DOB2(mdout1_1_20), 
        .DOB1(mdout1_1_19), .DOB0(mdout1_1_18))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7 (.DIA8(Data[35]), 
        .DIA7(Data[34]), .DIA6(Data[33]), .DIA5(Data[32]), .DIA4(Data[31]), 
        .DIA3(Data[30]), .DIA2(Data[29]), .DIA1(Data[28]), .DIA0(Data[27]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_35), .DOB7(mdout1_1_34), .DOB6(mdout1_1_33), 
        .DOB5(mdout1_1_32), .DOB4(mdout1_1_31), .DOB3(mdout1_1_30), .DOB2(mdout1_1_29), 
        .DOB1(mdout1_1_28), .DOB0(mdout1_1_27))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6 (.DIA8(Data[44]), 
        .DIA7(Data[43]), .DIA6(Data[42]), .DIA5(Data[41]), .DIA4(Data[40]), 
        .DIA3(Data[39]), .DIA2(Data[38]), .DIA1(Data[37]), .DIA0(Data[36]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_44), .DOB7(mdout1_1_43), .DOB6(mdout1_1_42), 
        .DOB5(mdout1_1_41), .DOB4(mdout1_1_40), .DOB3(mdout1_1_39), .DOB2(mdout1_1_38), 
        .DOB1(mdout1_1_37), .DOB0(mdout1_1_36))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5 (.DIA8(Data[53]), 
        .DIA7(Data[52]), .DIA6(Data[51]), .DIA5(Data[50]), .DIA4(Data[49]), 
        .DIA3(Data[48]), .DIA2(Data[47]), .DIA1(Data[46]), .DIA0(Data[45]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_53), .DOB7(mdout1_1_52), .DOB6(mdout1_1_51), 
        .DOB5(mdout1_1_50), .DOB4(mdout1_1_49), .DOB3(mdout1_1_48), .DOB2(mdout1_1_47), 
        .DOB1(mdout1_1_46), .DOB0(mdout1_1_45))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4 (.DIA8(Data[62]), 
        .DIA7(Data[61]), .DIA6(Data[60]), .DIA5(Data[59]), .DIA4(Data[58]), 
        .DIA3(Data[57]), .DIA2(Data[56]), .DIA1(Data[55]), .DIA0(Data[54]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_62), .DOB7(mdout1_1_61), .DOB6(mdout1_1_60), 
        .DOB5(mdout1_1_59), .DOB4(mdout1_1_58), .DOB3(mdout1_1_57), .DOB2(mdout1_1_56), 
        .DOB1(mdout1_1_55), .DOB0(mdout1_1_54))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3 (.DIA8(Data[71]), 
        .DIA7(Data[70]), .DIA6(Data[69]), .DIA5(Data[68]), .DIA4(Data[67]), 
        .DIA3(Data[66]), .DIA2(Data[65]), .DIA1(Data[64]), .DIA0(Data[63]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_71), .DOB7(mdout1_1_70), .DOB6(mdout1_1_69), 
        .DOB5(mdout1_1_68), .DOB4(mdout1_1_67), .DOB3(mdout1_1_66), .DOB2(mdout1_1_65), 
        .DOB1(mdout1_1_64), .DOB0(mdout1_1_63))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2 (.DIA8(Data[80]), 
        .DIA7(Data[79]), .DIA6(Data[78]), .DIA5(Data[77]), .DIA4(Data[76]), 
        .DIA3(Data[75]), .DIA2(Data[74]), .DIA1(Data[73]), .DIA0(Data[72]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_80), .DOB7(mdout1_1_79), .DOB6(mdout1_1_78), 
        .DOB5(mdout1_1_77), .DOB4(mdout1_1_76), .DOB3(mdout1_1_75), .DOB2(mdout1_1_74), 
        .DOB1(mdout1_1_73), .DOB0(mdout1_1_72))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1 (.DIA8(Data[89]), 
        .DIA7(Data[88]), .DIA6(Data[87]), .DIA5(Data[86]), .DIA4(Data[85]), 
        .DIA3(Data[84]), .DIA2(Data[83]), .DIA1(Data[82]), .DIA0(Data[81]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(mdout1_1_89), .DOB7(mdout1_1_88), .DOB6(mdout1_1_87), 
        .DOB5(mdout1_1_86), .DOB4(mdout1_1_85), .DOB3(mdout1_1_84), .DOB2(mdout1_1_83), 
        .DOB1(mdout1_1_82), .DOB0(mdout1_1_81))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.INIT_DATA = "STATIC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.ASYNC_RESET_RELEASE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.CSDECODE_B = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.CSDECODE_A = "0b001" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.WRITEMODE_B = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.WRITEMODE_A = "NORMAL" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.GSR = "ENABLED" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.RESETMODE = "ASYNC" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.REGMODE_B = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.REGMODE_A = "OUTREG" ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.DATA_WIDTH_B = 9 ;
    defparam pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0.DATA_WIDTH_A = 9 ;
    DP8KC pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0 (.DIA8(scuba_vlo), 
        .DIA7(scuba_vlo), .DIA6(scuba_vlo), .DIA5(scuba_vlo), .DIA4(scuba_vlo), 
        .DIA3(scuba_vlo), .DIA2(scuba_vlo), .DIA1(scuba_vlo), .DIA0(Data[90]), 
        .ADA12(WrAddress[9]), .ADA11(WrAddress[8]), .ADA10(WrAddress[7]), 
        .ADA9(WrAddress[6]), .ADA8(WrAddress[5]), .ADA7(WrAddress[4]), .ADA6(WrAddress[3]), 
        .ADA5(WrAddress[2]), .ADA4(WrAddress[1]), .ADA3(WrAddress[0]), .ADA2(scuba_vlo), 
        .ADA1(scuba_vlo), .ADA0(scuba_vhi), .CEA(WrClockEn), .OCEA(WrClockEn), 
        .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo), .CSA0(WrAddress[10]), 
        .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo), .DIB6(scuba_vlo), 
        .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo), .DIB2(scuba_vlo), 
        .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(RdAddress[9]), .ADB11(RdAddress[8]), 
        .ADB10(RdAddress[7]), .ADB9(RdAddress[6]), .ADB8(RdAddress[5]), 
        .ADB7(RdAddress[4]), .ADB6(RdAddress[3]), .ADB5(RdAddress[2]), .ADB4(RdAddress[1]), 
        .ADB3(RdAddress[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo), 
        .CEB(RdClockEn), .OCEB(RdClockEn), .CLKB(RdClock), .WEB(scuba_vlo), 
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(RdAddress[10]), .RSTB(Reset), 
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(), .DOA2(), .DOA1(), 
        .DOA0(), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(), .DOB3(), .DOB2(), 
        .DOB1(), .DOB0(mdout1_1_90))
             /* synthesis MEM_LPC_FILE="pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B" */
             /* synthesis MEM_INIT_FILE="" */;

    FD1P3DX FF_1 (.D(RdAddress[10]), .SP(RdClockEn), .CK(RdClock), .CD(scuba_vlo), 
        .Q(raddr10_ff))
             /* synthesis GSR="ENABLED" */;

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    FD1P3DX FF_0 (.D(raddr10_ff), .SP(RdClockEn), .CK(RdClock), .CD(scuba_vlo), 
        .Q(raddr10_ff2))
             /* synthesis GSR="ENABLED" */;

    MUX21 mux_90 (.D0(mdout1_0_0), .D1(mdout1_1_0), .SD(raddr10_ff2), .Z(Q[0]));

    MUX21 mux_89 (.D0(mdout1_0_1), .D1(mdout1_1_1), .SD(raddr10_ff2), .Z(Q[1]));

    MUX21 mux_88 (.D0(mdout1_0_2), .D1(mdout1_1_2), .SD(raddr10_ff2), .Z(Q[2]));

    MUX21 mux_87 (.D0(mdout1_0_3), .D1(mdout1_1_3), .SD(raddr10_ff2), .Z(Q[3]));

    MUX21 mux_86 (.D0(mdout1_0_4), .D1(mdout1_1_4), .SD(raddr10_ff2), .Z(Q[4]));

    MUX21 mux_85 (.D0(mdout1_0_5), .D1(mdout1_1_5), .SD(raddr10_ff2), .Z(Q[5]));

    MUX21 mux_84 (.D0(mdout1_0_6), .D1(mdout1_1_6), .SD(raddr10_ff2), .Z(Q[6]));

    MUX21 mux_83 (.D0(mdout1_0_7), .D1(mdout1_1_7), .SD(raddr10_ff2), .Z(Q[7]));

    MUX21 mux_82 (.D0(mdout1_0_8), .D1(mdout1_1_8), .SD(raddr10_ff2), .Z(Q[8]));

    MUX21 mux_81 (.D0(mdout1_0_9), .D1(mdout1_1_9), .SD(raddr10_ff2), .Z(Q[9]));

    MUX21 mux_80 (.D0(mdout1_0_10), .D1(mdout1_1_10), .SD(raddr10_ff2), 
        .Z(Q[10]));

    MUX21 mux_79 (.D0(mdout1_0_11), .D1(mdout1_1_11), .SD(raddr10_ff2), 
        .Z(Q[11]));

    MUX21 mux_78 (.D0(mdout1_0_12), .D1(mdout1_1_12), .SD(raddr10_ff2), 
        .Z(Q[12]));

    MUX21 mux_77 (.D0(mdout1_0_13), .D1(mdout1_1_13), .SD(raddr10_ff2), 
        .Z(Q[13]));

    MUX21 mux_76 (.D0(mdout1_0_14), .D1(mdout1_1_14), .SD(raddr10_ff2), 
        .Z(Q[14]));

    MUX21 mux_75 (.D0(mdout1_0_15), .D1(mdout1_1_15), .SD(raddr10_ff2), 
        .Z(Q[15]));

    MUX21 mux_74 (.D0(mdout1_0_16), .D1(mdout1_1_16), .SD(raddr10_ff2), 
        .Z(Q[16]));

    MUX21 mux_73 (.D0(mdout1_0_17), .D1(mdout1_1_17), .SD(raddr10_ff2), 
        .Z(Q[17]));

    MUX21 mux_72 (.D0(mdout1_0_18), .D1(mdout1_1_18), .SD(raddr10_ff2), 
        .Z(Q[18]));

    MUX21 mux_71 (.D0(mdout1_0_19), .D1(mdout1_1_19), .SD(raddr10_ff2), 
        .Z(Q[19]));

    MUX21 mux_70 (.D0(mdout1_0_20), .D1(mdout1_1_20), .SD(raddr10_ff2), 
        .Z(Q[20]));

    MUX21 mux_69 (.D0(mdout1_0_21), .D1(mdout1_1_21), .SD(raddr10_ff2), 
        .Z(Q[21]));

    MUX21 mux_68 (.D0(mdout1_0_22), .D1(mdout1_1_22), .SD(raddr10_ff2), 
        .Z(Q[22]));

    MUX21 mux_67 (.D0(mdout1_0_23), .D1(mdout1_1_23), .SD(raddr10_ff2), 
        .Z(Q[23]));

    MUX21 mux_66 (.D0(mdout1_0_24), .D1(mdout1_1_24), .SD(raddr10_ff2), 
        .Z(Q[24]));

    MUX21 mux_65 (.D0(mdout1_0_25), .D1(mdout1_1_25), .SD(raddr10_ff2), 
        .Z(Q[25]));

    MUX21 mux_64 (.D0(mdout1_0_26), .D1(mdout1_1_26), .SD(raddr10_ff2), 
        .Z(Q[26]));

    MUX21 mux_63 (.D0(mdout1_0_27), .D1(mdout1_1_27), .SD(raddr10_ff2), 
        .Z(Q[27]));

    MUX21 mux_62 (.D0(mdout1_0_28), .D1(mdout1_1_28), .SD(raddr10_ff2), 
        .Z(Q[28]));

    MUX21 mux_61 (.D0(mdout1_0_29), .D1(mdout1_1_29), .SD(raddr10_ff2), 
        .Z(Q[29]));

    MUX21 mux_60 (.D0(mdout1_0_30), .D1(mdout1_1_30), .SD(raddr10_ff2), 
        .Z(Q[30]));

    MUX21 mux_59 (.D0(mdout1_0_31), .D1(mdout1_1_31), .SD(raddr10_ff2), 
        .Z(Q[31]));

    MUX21 mux_58 (.D0(mdout1_0_32), .D1(mdout1_1_32), .SD(raddr10_ff2), 
        .Z(Q[32]));

    MUX21 mux_57 (.D0(mdout1_0_33), .D1(mdout1_1_33), .SD(raddr10_ff2), 
        .Z(Q[33]));

    MUX21 mux_56 (.D0(mdout1_0_34), .D1(mdout1_1_34), .SD(raddr10_ff2), 
        .Z(Q[34]));

    MUX21 mux_55 (.D0(mdout1_0_35), .D1(mdout1_1_35), .SD(raddr10_ff2), 
        .Z(Q[35]));

    MUX21 mux_54 (.D0(mdout1_0_36), .D1(mdout1_1_36), .SD(raddr10_ff2), 
        .Z(Q[36]));

    MUX21 mux_53 (.D0(mdout1_0_37), .D1(mdout1_1_37), .SD(raddr10_ff2), 
        .Z(Q[37]));

    MUX21 mux_52 (.D0(mdout1_0_38), .D1(mdout1_1_38), .SD(raddr10_ff2), 
        .Z(Q[38]));

    MUX21 mux_51 (.D0(mdout1_0_39), .D1(mdout1_1_39), .SD(raddr10_ff2), 
        .Z(Q[39]));

    MUX21 mux_50 (.D0(mdout1_0_40), .D1(mdout1_1_40), .SD(raddr10_ff2), 
        .Z(Q[40]));

    MUX21 mux_49 (.D0(mdout1_0_41), .D1(mdout1_1_41), .SD(raddr10_ff2), 
        .Z(Q[41]));

    MUX21 mux_48 (.D0(mdout1_0_42), .D1(mdout1_1_42), .SD(raddr10_ff2), 
        .Z(Q[42]));

    MUX21 mux_47 (.D0(mdout1_0_43), .D1(mdout1_1_43), .SD(raddr10_ff2), 
        .Z(Q[43]));

    MUX21 mux_46 (.D0(mdout1_0_44), .D1(mdout1_1_44), .SD(raddr10_ff2), 
        .Z(Q[44]));

    MUX21 mux_45 (.D0(mdout1_0_45), .D1(mdout1_1_45), .SD(raddr10_ff2), 
        .Z(Q[45]));

    MUX21 mux_44 (.D0(mdout1_0_46), .D1(mdout1_1_46), .SD(raddr10_ff2), 
        .Z(Q[46]));

    MUX21 mux_43 (.D0(mdout1_0_47), .D1(mdout1_1_47), .SD(raddr10_ff2), 
        .Z(Q[47]));

    MUX21 mux_42 (.D0(mdout1_0_48), .D1(mdout1_1_48), .SD(raddr10_ff2), 
        .Z(Q[48]));

    MUX21 mux_41 (.D0(mdout1_0_49), .D1(mdout1_1_49), .SD(raddr10_ff2), 
        .Z(Q[49]));

    MUX21 mux_40 (.D0(mdout1_0_50), .D1(mdout1_1_50), .SD(raddr10_ff2), 
        .Z(Q[50]));

    MUX21 mux_39 (.D0(mdout1_0_51), .D1(mdout1_1_51), .SD(raddr10_ff2), 
        .Z(Q[51]));

    MUX21 mux_38 (.D0(mdout1_0_52), .D1(mdout1_1_52), .SD(raddr10_ff2), 
        .Z(Q[52]));

    MUX21 mux_37 (.D0(mdout1_0_53), .D1(mdout1_1_53), .SD(raddr10_ff2), 
        .Z(Q[53]));

    MUX21 mux_36 (.D0(mdout1_0_54), .D1(mdout1_1_54), .SD(raddr10_ff2), 
        .Z(Q[54]));

    MUX21 mux_35 (.D0(mdout1_0_55), .D1(mdout1_1_55), .SD(raddr10_ff2), 
        .Z(Q[55]));

    MUX21 mux_34 (.D0(mdout1_0_56), .D1(mdout1_1_56), .SD(raddr10_ff2), 
        .Z(Q[56]));

    MUX21 mux_33 (.D0(mdout1_0_57), .D1(mdout1_1_57), .SD(raddr10_ff2), 
        .Z(Q[57]));

    MUX21 mux_32 (.D0(mdout1_0_58), .D1(mdout1_1_58), .SD(raddr10_ff2), 
        .Z(Q[58]));

    MUX21 mux_31 (.D0(mdout1_0_59), .D1(mdout1_1_59), .SD(raddr10_ff2), 
        .Z(Q[59]));

    MUX21 mux_30 (.D0(mdout1_0_60), .D1(mdout1_1_60), .SD(raddr10_ff2), 
        .Z(Q[60]));

    MUX21 mux_29 (.D0(mdout1_0_61), .D1(mdout1_1_61), .SD(raddr10_ff2), 
        .Z(Q[61]));

    MUX21 mux_28 (.D0(mdout1_0_62), .D1(mdout1_1_62), .SD(raddr10_ff2), 
        .Z(Q[62]));

    MUX21 mux_27 (.D0(mdout1_0_63), .D1(mdout1_1_63), .SD(raddr10_ff2), 
        .Z(Q[63]));

    MUX21 mux_26 (.D0(mdout1_0_64), .D1(mdout1_1_64), .SD(raddr10_ff2), 
        .Z(Q[64]));

    MUX21 mux_25 (.D0(mdout1_0_65), .D1(mdout1_1_65), .SD(raddr10_ff2), 
        .Z(Q[65]));

    MUX21 mux_24 (.D0(mdout1_0_66), .D1(mdout1_1_66), .SD(raddr10_ff2), 
        .Z(Q[66]));

    MUX21 mux_23 (.D0(mdout1_0_67), .D1(mdout1_1_67), .SD(raddr10_ff2), 
        .Z(Q[67]));

    MUX21 mux_22 (.D0(mdout1_0_68), .D1(mdout1_1_68), .SD(raddr10_ff2), 
        .Z(Q[68]));

    MUX21 mux_21 (.D0(mdout1_0_69), .D1(mdout1_1_69), .SD(raddr10_ff2), 
        .Z(Q[69]));

    MUX21 mux_20 (.D0(mdout1_0_70), .D1(mdout1_1_70), .SD(raddr10_ff2), 
        .Z(Q[70]));

    MUX21 mux_19 (.D0(mdout1_0_71), .D1(mdout1_1_71), .SD(raddr10_ff2), 
        .Z(Q[71]));

    MUX21 mux_18 (.D0(mdout1_0_72), .D1(mdout1_1_72), .SD(raddr10_ff2), 
        .Z(Q[72]));

    MUX21 mux_17 (.D0(mdout1_0_73), .D1(mdout1_1_73), .SD(raddr10_ff2), 
        .Z(Q[73]));

    MUX21 mux_16 (.D0(mdout1_0_74), .D1(mdout1_1_74), .SD(raddr10_ff2), 
        .Z(Q[74]));

    MUX21 mux_15 (.D0(mdout1_0_75), .D1(mdout1_1_75), .SD(raddr10_ff2), 
        .Z(Q[75]));

    MUX21 mux_14 (.D0(mdout1_0_76), .D1(mdout1_1_76), .SD(raddr10_ff2), 
        .Z(Q[76]));

    MUX21 mux_13 (.D0(mdout1_0_77), .D1(mdout1_1_77), .SD(raddr10_ff2), 
        .Z(Q[77]));

    MUX21 mux_12 (.D0(mdout1_0_78), .D1(mdout1_1_78), .SD(raddr10_ff2), 
        .Z(Q[78]));

    MUX21 mux_11 (.D0(mdout1_0_79), .D1(mdout1_1_79), .SD(raddr10_ff2), 
        .Z(Q[79]));

    MUX21 mux_10 (.D0(mdout1_0_80), .D1(mdout1_1_80), .SD(raddr10_ff2), 
        .Z(Q[80]));

    MUX21 mux_9 (.D0(mdout1_0_81), .D1(mdout1_1_81), .SD(raddr10_ff2), .Z(Q[81]));

    MUX21 mux_8 (.D0(mdout1_0_82), .D1(mdout1_1_82), .SD(raddr10_ff2), .Z(Q[82]));

    MUX21 mux_7 (.D0(mdout1_0_83), .D1(mdout1_1_83), .SD(raddr10_ff2), .Z(Q[83]));

    MUX21 mux_6 (.D0(mdout1_0_84), .D1(mdout1_1_84), .SD(raddr10_ff2), .Z(Q[84]));

    MUX21 mux_5 (.D0(mdout1_0_85), .D1(mdout1_1_85), .SD(raddr10_ff2), .Z(Q[85]));

    MUX21 mux_4 (.D0(mdout1_0_86), .D1(mdout1_1_86), .SD(raddr10_ff2), .Z(Q[86]));

    MUX21 mux_3 (.D0(mdout1_0_87), .D1(mdout1_1_87), .SD(raddr10_ff2), .Z(Q[87]));

    MUX21 mux_2 (.D0(mdout1_0_88), .D1(mdout1_1_88), .SD(raddr10_ff2), .Z(Q[88]));

    MUX21 mux_1 (.D0(mdout1_0_89), .D1(mdout1_1_89), .SD(raddr10_ff2), .Z(Q[89]));

    MUX21 mux_0 (.D0(mdout1_0_90), .D1(mdout1_1_90), .SD(raddr10_ff2), .Z(Q[90]));



    // exemplar begin
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_0_21 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_1_20 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_2_19 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_3_18 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_4_17 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_5_16 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_6_15 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_7_14 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_8_13 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_9_12 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_0_10_11 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_0_10 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_1_9 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_2_8 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_3_7 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_4_6 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_5_5 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_6_4 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_7_3 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_8_2 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_9_1 MEM_INIT_FILE 
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0 MEM_LPC_FILE pmi_ram_dpXbnonesadr911120489111204811f45a5e__PMIP__2048__91__91B
    // exemplar attribute pmi_ram_dpXbnonesadr911120489111204811f45a5e_1_10_0 MEM_INIT_FILE 
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar end

endmodule
